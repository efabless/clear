magic
tech sky130A
magscale 1 2
timestamp 1656943463
<< viali >>
rect 1961 20553 1995 20587
rect 21005 20553 21039 20587
rect 2145 20417 2179 20451
rect 14105 20417 14139 20451
rect 17785 20417 17819 20451
rect 20269 20417 20303 20451
rect 20821 20417 20855 20451
rect 7849 20349 7883 20383
rect 14289 20349 14323 20383
rect 17141 20349 17175 20383
rect 17877 20349 17911 20383
rect 18061 20349 18095 20383
rect 2513 20213 2547 20247
rect 12357 20213 12391 20247
rect 17417 20213 17451 20247
rect 18429 20213 18463 20247
rect 19901 20213 19935 20247
rect 20453 20213 20487 20247
rect 2513 20009 2547 20043
rect 13737 20009 13771 20043
rect 14105 20009 14139 20043
rect 20913 20009 20947 20043
rect 12725 19941 12759 19975
rect 3985 19873 4019 19907
rect 7665 19873 7699 19907
rect 10517 19873 10551 19907
rect 11897 19873 11931 19907
rect 14749 19873 14783 19907
rect 16681 19873 16715 19907
rect 17325 19873 17359 19907
rect 18245 19873 18279 19907
rect 2145 19805 2179 19839
rect 2697 19805 2731 19839
rect 2973 19805 3007 19839
rect 4261 19805 4295 19839
rect 7849 19805 7883 19839
rect 11805 19805 11839 19839
rect 12541 19805 12575 19839
rect 13093 19805 13127 19839
rect 14565 19805 14599 19839
rect 15117 19805 15151 19839
rect 16497 19805 16531 19839
rect 19257 19805 19291 19839
rect 19533 19805 19567 19839
rect 19993 19805 20027 19839
rect 20729 19805 20763 19839
rect 21281 19805 21315 19839
rect 10333 19737 10367 19771
rect 14473 19737 14507 19771
rect 15393 19737 15427 19771
rect 1961 19669 1995 19703
rect 7113 19669 7147 19703
rect 7757 19669 7791 19703
rect 8217 19669 8251 19703
rect 9965 19669 9999 19703
rect 10425 19669 10459 19703
rect 11069 19669 11103 19703
rect 11345 19669 11379 19703
rect 11713 19669 11747 19703
rect 13277 19669 13311 19703
rect 16129 19669 16163 19703
rect 16589 19669 16623 19703
rect 17509 19669 17543 19703
rect 17601 19669 17635 19703
rect 17969 19669 18003 19703
rect 18705 19669 18739 19703
rect 20177 19669 20211 19703
rect 2513 19465 2547 19499
rect 4721 19465 4755 19499
rect 7941 19465 7975 19499
rect 10425 19465 10459 19499
rect 11805 19465 11839 19499
rect 14841 19465 14875 19499
rect 16037 19465 16071 19499
rect 17141 19465 17175 19499
rect 17417 19465 17451 19499
rect 17785 19465 17819 19499
rect 14381 19397 14415 19431
rect 1593 19329 1627 19363
rect 2145 19329 2179 19363
rect 2697 19329 2731 19363
rect 5089 19329 5123 19363
rect 5181 19329 5215 19363
rect 10057 19329 10091 19363
rect 14473 19329 14507 19363
rect 20729 19329 20763 19363
rect 2973 19261 3007 19295
rect 5365 19261 5399 19295
rect 6469 19261 6503 19295
rect 8033 19261 8067 19295
rect 8217 19261 8251 19295
rect 9413 19261 9447 19295
rect 9873 19261 9907 19295
rect 9965 19261 9999 19295
rect 10701 19261 10735 19295
rect 12357 19261 12391 19295
rect 14289 19261 14323 19295
rect 17877 19261 17911 19295
rect 17969 19261 18003 19295
rect 1961 19193 1995 19227
rect 5825 19193 5859 19227
rect 16681 19193 16715 19227
rect 6745 19125 6779 19159
rect 7573 19125 7607 19159
rect 15393 19125 15427 19159
rect 20913 19125 20947 19159
rect 5273 18921 5307 18955
rect 14565 18921 14599 18955
rect 16589 18921 16623 18955
rect 18521 18921 18555 18955
rect 3801 18853 3835 18887
rect 19993 18853 20027 18887
rect 4445 18785 4479 18819
rect 5917 18785 5951 18819
rect 8953 18785 8987 18819
rect 11989 18785 12023 18819
rect 12633 18785 12667 18819
rect 15117 18785 15151 18819
rect 16129 18785 16163 18819
rect 17233 18785 17267 18819
rect 19349 18785 19383 18819
rect 19533 18785 19567 18819
rect 2145 18717 2179 18751
rect 3065 18717 3099 18751
rect 3341 18717 3375 18751
rect 4169 18717 4203 18751
rect 7941 18717 7975 18751
rect 11805 18717 11839 18751
rect 15945 18717 15979 18751
rect 17049 18717 17083 18751
rect 20821 18717 20855 18751
rect 5641 18649 5675 18683
rect 6285 18649 6319 18683
rect 7113 18649 7147 18683
rect 12725 18649 12759 18683
rect 14933 18649 14967 18683
rect 16957 18649 16991 18683
rect 18061 18649 18095 18683
rect 1961 18581 1995 18615
rect 2605 18581 2639 18615
rect 4261 18581 4295 18615
rect 5733 18581 5767 18615
rect 6745 18581 6779 18615
rect 7573 18581 7607 18615
rect 9505 18581 9539 18615
rect 9873 18581 9907 18615
rect 11069 18581 11103 18615
rect 11437 18581 11471 18615
rect 11897 18581 11931 18615
rect 12817 18581 12851 18615
rect 13185 18581 13219 18615
rect 15025 18581 15059 18615
rect 15577 18581 15611 18615
rect 16037 18581 16071 18615
rect 17601 18581 17635 18615
rect 19625 18581 19659 18615
rect 20361 18581 20395 18615
rect 21005 18581 21039 18615
rect 3617 18377 3651 18411
rect 4261 18377 4295 18411
rect 5733 18377 5767 18411
rect 7941 18377 7975 18411
rect 8309 18377 8343 18411
rect 10149 18377 10183 18411
rect 12357 18377 12391 18411
rect 13829 18377 13863 18411
rect 15393 18377 15427 18411
rect 18061 18377 18095 18411
rect 18153 18377 18187 18411
rect 7665 18309 7699 18343
rect 19165 18309 19199 18343
rect 1593 18241 1627 18275
rect 2145 18241 2179 18275
rect 3249 18241 3283 18275
rect 4997 18241 5031 18275
rect 5641 18241 5675 18275
rect 8401 18241 8435 18275
rect 9321 18241 9355 18275
rect 9965 18241 9999 18275
rect 11161 18241 11195 18275
rect 11989 18241 12023 18275
rect 12633 18241 12667 18275
rect 13645 18241 13679 18275
rect 14197 18241 14231 18275
rect 15301 18241 15335 18275
rect 20269 18241 20303 18275
rect 20821 18241 20855 18275
rect 2973 18173 3007 18207
rect 3157 18173 3191 18207
rect 3985 18173 4019 18207
rect 4169 18173 4203 18207
rect 5917 18173 5951 18207
rect 8493 18173 8527 18207
rect 9413 18173 9447 18207
rect 9505 18173 9539 18207
rect 11713 18173 11747 18207
rect 11897 18173 11931 18207
rect 13185 18173 13219 18207
rect 15577 18173 15611 18207
rect 17969 18173 18003 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 5273 18105 5307 18139
rect 16773 18105 16807 18139
rect 1961 18037 1995 18071
rect 2421 18037 2455 18071
rect 4629 18037 4663 18071
rect 6653 18037 6687 18071
rect 7297 18037 7331 18071
rect 8953 18037 8987 18071
rect 10609 18037 10643 18071
rect 14933 18037 14967 18071
rect 16221 18037 16255 18071
rect 17233 18037 17267 18071
rect 18521 18037 18555 18071
rect 18797 18037 18831 18071
rect 19809 18037 19843 18071
rect 20453 18037 20487 18071
rect 21005 18037 21039 18071
rect 1961 17833 1995 17867
rect 2605 17833 2639 17867
rect 5641 17833 5675 17867
rect 9597 17833 9631 17867
rect 16129 17833 16163 17867
rect 16589 17833 16623 17867
rect 19257 17833 19291 17867
rect 21281 17833 21315 17867
rect 11529 17765 11563 17799
rect 17601 17765 17635 17799
rect 3801 17697 3835 17731
rect 4813 17697 4847 17731
rect 6285 17697 6319 17731
rect 6929 17697 6963 17731
rect 7941 17697 7975 17731
rect 10241 17697 10275 17731
rect 12081 17697 12115 17731
rect 13001 17697 13035 17731
rect 15577 17697 15611 17731
rect 18245 17697 18279 17731
rect 19809 17697 19843 17731
rect 20821 17697 20855 17731
rect 2145 17629 2179 17663
rect 2789 17629 2823 17663
rect 4261 17629 4295 17663
rect 16405 17629 16439 17663
rect 16957 17629 16991 17663
rect 17969 17629 18003 17663
rect 19625 17629 19659 17663
rect 4905 17561 4939 17595
rect 8033 17561 8067 17595
rect 8125 17561 8159 17595
rect 8953 17561 8987 17595
rect 10057 17561 10091 17595
rect 11161 17561 11195 17595
rect 11897 17561 11931 17595
rect 12541 17561 12575 17595
rect 1593 17493 1627 17527
rect 3065 17493 3099 17527
rect 4997 17493 5031 17527
rect 5365 17493 5399 17527
rect 6009 17493 6043 17527
rect 6101 17493 6135 17527
rect 7021 17493 7055 17527
rect 7113 17493 7147 17527
rect 7481 17493 7515 17527
rect 8493 17493 8527 17527
rect 9965 17493 9999 17527
rect 10793 17493 10827 17527
rect 11989 17493 12023 17527
rect 15025 17493 15059 17527
rect 15669 17493 15703 17527
rect 15761 17493 15795 17527
rect 18061 17493 18095 17527
rect 18613 17493 18647 17527
rect 19717 17493 19751 17527
rect 20269 17493 20303 17527
rect 20637 17493 20671 17527
rect 20729 17493 20763 17527
rect 1501 17289 1535 17323
rect 4445 17289 4479 17323
rect 5181 17289 5215 17323
rect 6837 17289 6871 17323
rect 8401 17289 8435 17323
rect 8493 17289 8527 17323
rect 9045 17289 9079 17323
rect 10701 17289 10735 17323
rect 14289 17289 14323 17323
rect 14749 17289 14783 17323
rect 20821 17289 20855 17323
rect 3985 17221 4019 17255
rect 5089 17221 5123 17255
rect 19809 17221 19843 17255
rect 20729 17221 20763 17255
rect 1685 17153 1719 17187
rect 1961 17153 1995 17187
rect 2973 17153 3007 17187
rect 3433 17153 3467 17187
rect 4077 17153 4111 17187
rect 6929 17153 6963 17187
rect 7573 17153 7607 17187
rect 9413 17153 9447 17187
rect 10793 17153 10827 17187
rect 11989 17153 12023 17187
rect 12633 17153 12667 17187
rect 14381 17153 14415 17187
rect 15025 17153 15059 17187
rect 16681 17153 16715 17187
rect 17233 17153 17267 17187
rect 20085 17153 20119 17187
rect 3893 17085 3927 17119
rect 5365 17085 5399 17119
rect 6745 17085 6779 17119
rect 8677 17085 8711 17119
rect 9505 17085 9539 17119
rect 9597 17085 9631 17119
rect 10609 17085 10643 17119
rect 11805 17085 11839 17119
rect 11897 17085 11931 17119
rect 14197 17085 14231 17119
rect 18061 17085 18095 17119
rect 20913 17085 20947 17119
rect 16865 17017 16899 17051
rect 2145 16949 2179 16983
rect 2789 16949 2823 16983
rect 4721 16949 4755 16983
rect 5917 16949 5951 16983
rect 7297 16949 7331 16983
rect 8033 16949 8067 16983
rect 10057 16949 10091 16983
rect 11161 16949 11195 16983
rect 12357 16949 12391 16983
rect 13645 16949 13679 16983
rect 17601 16949 17635 16983
rect 18521 16949 18555 16983
rect 20361 16949 20395 16983
rect 3341 16745 3375 16779
rect 7205 16745 7239 16779
rect 9137 16745 9171 16779
rect 16221 16745 16255 16779
rect 19993 16745 20027 16779
rect 4537 16677 4571 16711
rect 6193 16677 6227 16711
rect 8585 16677 8619 16711
rect 1961 16609 1995 16643
rect 3985 16609 4019 16643
rect 6561 16609 6595 16643
rect 9505 16609 9539 16643
rect 10057 16609 10091 16643
rect 11069 16609 11103 16643
rect 11897 16609 11931 16643
rect 12817 16609 12851 16643
rect 12909 16609 12943 16643
rect 15853 16609 15887 16643
rect 16681 16609 16715 16643
rect 16865 16609 16899 16643
rect 17785 16609 17819 16643
rect 20453 16609 20487 16643
rect 20545 16609 20579 16643
rect 2237 16541 2271 16575
rect 2973 16541 3007 16575
rect 8125 16541 8159 16575
rect 10241 16541 10275 16575
rect 11253 16541 11287 16575
rect 13001 16541 13035 16575
rect 17601 16541 17635 16575
rect 18797 16541 18831 16575
rect 21005 16541 21039 16575
rect 2697 16473 2731 16507
rect 4077 16473 4111 16507
rect 5825 16473 5859 16507
rect 7757 16473 7791 16507
rect 17693 16473 17727 16507
rect 18521 16473 18555 16507
rect 4169 16405 4203 16439
rect 4905 16405 4939 16439
rect 5273 16405 5307 16439
rect 6929 16405 6963 16439
rect 10149 16405 10183 16439
rect 10609 16405 10643 16439
rect 11161 16405 11195 16439
rect 11621 16405 11655 16439
rect 13369 16405 13403 16439
rect 16589 16405 16623 16439
rect 17233 16405 17267 16439
rect 20361 16405 20395 16439
rect 21189 16405 21223 16439
rect 2421 16201 2455 16235
rect 5089 16201 5123 16235
rect 5457 16201 5491 16235
rect 6561 16201 6595 16235
rect 7573 16201 7607 16235
rect 11529 16201 11563 16235
rect 14197 16201 14231 16235
rect 14565 16201 14599 16235
rect 16773 16201 16807 16235
rect 17693 16201 17727 16235
rect 18337 16201 18371 16235
rect 18797 16201 18831 16235
rect 7021 16133 7055 16167
rect 10250 16133 10284 16167
rect 20637 16133 20671 16167
rect 2053 16065 2087 16099
rect 2605 16065 2639 16099
rect 4445 16065 4479 16099
rect 5549 16065 5583 16099
rect 6929 16065 6963 16099
rect 7941 16065 7975 16099
rect 18705 16065 18739 16099
rect 20361 16065 20395 16099
rect 21097 16065 21131 16099
rect 4537 15997 4571 16031
rect 4721 15997 4755 16031
rect 5733 15997 5767 16031
rect 7113 15997 7147 16031
rect 8033 15997 8067 16031
rect 8217 15997 8251 16031
rect 10517 15997 10551 16031
rect 14013 15997 14047 16031
rect 14105 15997 14139 16031
rect 17509 15997 17543 16031
rect 17601 15997 17635 16031
rect 18981 15997 19015 16031
rect 19993 15997 20027 16031
rect 2973 15929 3007 15963
rect 18061 15929 18095 15963
rect 21281 15929 21315 15963
rect 1869 15861 1903 15895
rect 4077 15861 4111 15895
rect 8677 15861 8711 15895
rect 9137 15861 9171 15895
rect 10793 15861 10827 15895
rect 13461 15861 13495 15895
rect 14933 15861 14967 15895
rect 4445 15657 4479 15691
rect 8217 15657 8251 15691
rect 10609 15657 10643 15691
rect 13645 15657 13679 15691
rect 16957 15657 16991 15691
rect 19993 15657 20027 15691
rect 2329 15589 2363 15623
rect 6929 15589 6963 15623
rect 5089 15521 5123 15555
rect 6377 15521 6411 15555
rect 7665 15521 7699 15555
rect 18521 15521 18555 15555
rect 2513 15453 2547 15487
rect 3341 15453 3375 15487
rect 6561 15453 6595 15487
rect 9229 15453 9263 15487
rect 10885 15453 10919 15487
rect 16589 15453 16623 15487
rect 20729 15453 20763 15487
rect 4813 15385 4847 15419
rect 5457 15385 5491 15419
rect 6469 15385 6503 15419
rect 8493 15385 8527 15419
rect 9474 15385 9508 15419
rect 16344 15385 16378 15419
rect 20361 15385 20395 15419
rect 2973 15317 3007 15351
rect 4169 15317 4203 15351
rect 4905 15317 4939 15351
rect 7757 15317 7791 15351
rect 7849 15317 7883 15351
rect 15209 15317 15243 15351
rect 17325 15317 17359 15351
rect 19625 15317 19659 15351
rect 20913 15317 20947 15351
rect 21281 15317 21315 15351
rect 3893 15113 3927 15147
rect 14841 15113 14875 15147
rect 15945 15113 15979 15147
rect 7757 15045 7791 15079
rect 8309 15045 8343 15079
rect 20146 15045 20180 15079
rect 1869 14977 1903 15011
rect 2881 14977 2915 15011
rect 3157 14977 3191 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 7665 14977 7699 15011
rect 9689 14977 9723 15011
rect 9956 14977 9990 15011
rect 13461 14977 13495 15011
rect 13728 14977 13762 15011
rect 16681 14977 16715 15011
rect 16948 14977 16982 15011
rect 2145 14909 2179 14943
rect 5273 14909 5307 14943
rect 5917 14909 5951 14943
rect 7941 14909 7975 14943
rect 19901 14909 19935 14943
rect 6929 14841 6963 14875
rect 2697 14773 2731 14807
rect 3341 14773 3375 14807
rect 4261 14773 4295 14807
rect 4629 14773 4663 14807
rect 6653 14773 6687 14807
rect 7297 14773 7331 14807
rect 11069 14773 11103 14807
rect 11621 14773 11655 14807
rect 15209 14773 15243 14807
rect 15669 14773 15703 14807
rect 18061 14773 18095 14807
rect 18429 14773 18463 14807
rect 18889 14773 18923 14807
rect 19533 14773 19567 14807
rect 21281 14773 21315 14807
rect 5089 14569 5123 14603
rect 11897 14569 11931 14603
rect 14105 14569 14139 14603
rect 17141 14569 17175 14603
rect 17417 14569 17451 14603
rect 19257 14569 19291 14603
rect 21097 14569 21131 14603
rect 3433 14433 3467 14467
rect 4353 14433 4387 14467
rect 5733 14433 5767 14467
rect 7021 14433 7055 14467
rect 7205 14433 7239 14467
rect 10241 14433 10275 14467
rect 2145 14365 2179 14399
rect 2789 14365 2823 14399
rect 3065 14365 3099 14399
rect 7297 14365 7331 14399
rect 10508 14365 10542 14399
rect 13277 14365 13311 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 16028 14365 16062 14399
rect 18797 14365 18831 14399
rect 20637 14365 20671 14399
rect 20913 14365 20947 14399
rect 4261 14297 4295 14331
rect 5457 14297 5491 14331
rect 6469 14297 6503 14331
rect 13010 14297 13044 14331
rect 15218 14297 15252 14331
rect 18530 14297 18564 14331
rect 20370 14297 20404 14331
rect 1961 14229 1995 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 5549 14229 5583 14263
rect 6193 14229 6227 14263
rect 7665 14229 7699 14263
rect 11621 14229 11655 14263
rect 13645 14229 13679 14263
rect 3985 14025 4019 14059
rect 4445 14025 4479 14059
rect 5549 14025 5583 14059
rect 14289 14025 14323 14059
rect 15945 14025 15979 14059
rect 18981 14025 19015 14059
rect 19349 14025 19383 14059
rect 19901 14025 19935 14059
rect 3709 13957 3743 13991
rect 4353 13957 4387 13991
rect 6929 13957 6963 13991
rect 8125 13957 8159 13991
rect 14810 13957 14844 13991
rect 17868 13957 17902 13991
rect 1961 13889 1995 13923
rect 2421 13889 2455 13923
rect 2697 13889 2731 13923
rect 6837 13889 6871 13923
rect 8401 13889 8435 13923
rect 9229 13889 9263 13923
rect 9496 13889 9530 13923
rect 13165 13889 13199 13923
rect 17325 13889 17359 13923
rect 17601 13889 17635 13923
rect 21014 13889 21048 13923
rect 21281 13889 21315 13923
rect 4629 13821 4663 13855
rect 5825 13821 5859 13855
rect 7113 13821 7147 13855
rect 7757 13821 7791 13855
rect 10977 13821 11011 13855
rect 11713 13821 11747 13855
rect 12909 13821 12943 13855
rect 14565 13821 14599 13855
rect 16313 13821 16347 13855
rect 10609 13753 10643 13787
rect 1777 13685 1811 13719
rect 5089 13685 5123 13719
rect 6469 13685 6503 13719
rect 1685 13481 1719 13515
rect 3801 13481 3835 13515
rect 6469 13481 6503 13515
rect 10793 13481 10827 13515
rect 14473 13481 14507 13515
rect 17417 13481 17451 13515
rect 17693 13481 17727 13515
rect 21097 13481 21131 13515
rect 6193 13413 6227 13447
rect 2329 13345 2363 13379
rect 4445 13345 4479 13379
rect 5641 13345 5675 13379
rect 7021 13345 7055 13379
rect 8125 13345 8159 13379
rect 9413 13345 9447 13379
rect 5825 13277 5859 13311
rect 6929 13277 6963 13311
rect 16037 13277 16071 13311
rect 18797 13277 18831 13311
rect 20637 13277 20671 13311
rect 20913 13277 20947 13311
rect 4169 13209 4203 13243
rect 5181 13209 5215 13243
rect 5733 13209 5767 13243
rect 8953 13209 8987 13243
rect 9680 13209 9714 13243
rect 16304 13209 16338 13243
rect 20392 13209 20426 13243
rect 2053 13141 2087 13175
rect 2145 13141 2179 13175
rect 4261 13141 4295 13175
rect 6837 13141 6871 13175
rect 7481 13141 7515 13175
rect 7849 13141 7883 13175
rect 7941 13141 7975 13175
rect 8493 13141 8527 13175
rect 11161 13141 11195 13175
rect 19257 13141 19291 13175
rect 2421 12937 2455 12971
rect 5273 12937 5307 12971
rect 5733 12937 5767 12971
rect 7665 12937 7699 12971
rect 8677 12937 8711 12971
rect 9229 12937 9263 12971
rect 10977 12937 11011 12971
rect 11621 12937 11655 12971
rect 14105 12937 14139 12971
rect 15853 12937 15887 12971
rect 19257 12937 19291 12971
rect 20085 12937 20119 12971
rect 20545 12937 20579 12971
rect 4537 12869 4571 12903
rect 8309 12869 8343 12903
rect 10342 12869 10376 12903
rect 15240 12869 15274 12903
rect 19717 12869 19751 12903
rect 2053 12801 2087 12835
rect 3709 12801 3743 12835
rect 5641 12801 5675 12835
rect 7021 12801 7055 12835
rect 10609 12801 10643 12835
rect 13573 12801 13607 12835
rect 15485 12801 15519 12835
rect 17877 12801 17911 12835
rect 18144 12801 18178 12835
rect 20913 12801 20947 12835
rect 1777 12733 1811 12767
rect 1961 12733 1995 12767
rect 3525 12733 3559 12767
rect 3617 12733 3651 12767
rect 4905 12733 4939 12767
rect 5917 12733 5951 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 13829 12733 13863 12767
rect 21005 12733 21039 12767
rect 21097 12733 21131 12767
rect 4077 12597 4111 12631
rect 6561 12597 6595 12631
rect 7297 12597 7331 12631
rect 12449 12597 12483 12631
rect 3893 12393 3927 12427
rect 6929 12393 6963 12427
rect 12265 12393 12299 12427
rect 14473 12393 14507 12427
rect 17417 12393 17451 12427
rect 20085 12393 20119 12427
rect 21281 12393 21315 12427
rect 9229 12325 9263 12359
rect 2513 12257 2547 12291
rect 4445 12257 4479 12291
rect 6101 12257 6135 12291
rect 7573 12257 7607 12291
rect 10609 12257 10643 12291
rect 10885 12257 10919 12291
rect 20729 12257 20763 12291
rect 2329 12189 2363 12223
rect 7297 12189 7331 12223
rect 12633 12189 12667 12223
rect 14197 12189 14231 12223
rect 15669 12189 15703 12223
rect 20269 12189 20303 12223
rect 10342 12121 10376 12155
rect 11130 12121 11164 12155
rect 15936 12121 15970 12155
rect 17693 12121 17727 12155
rect 19349 12121 19383 12155
rect 20821 12121 20855 12155
rect 1501 12053 1535 12087
rect 1869 12053 1903 12087
rect 2237 12053 2271 12087
rect 2881 12053 2915 12087
rect 3249 12053 3283 12087
rect 4261 12053 4295 12087
rect 4353 12053 4387 12087
rect 4905 12053 4939 12087
rect 5273 12053 5307 12087
rect 6561 12053 6595 12087
rect 7389 12053 7423 12087
rect 8125 12053 8159 12087
rect 8493 12053 8527 12087
rect 17049 12053 17083 12087
rect 19625 12053 19659 12087
rect 20913 12053 20947 12087
rect 2053 11849 2087 11883
rect 2421 11849 2455 11883
rect 3065 11849 3099 11883
rect 3525 11849 3559 11883
rect 4261 11849 4295 11883
rect 5273 11849 5307 11883
rect 7205 11849 7239 11883
rect 9505 11849 9539 11883
rect 13185 11849 13219 11883
rect 19717 11849 19751 11883
rect 21189 11849 21223 11883
rect 4905 11781 4939 11815
rect 5641 11781 5675 11815
rect 7297 11781 7331 11815
rect 8677 11781 8711 11815
rect 12050 11781 12084 11815
rect 13553 11781 13587 11815
rect 15178 11781 15212 11815
rect 18236 11781 18270 11815
rect 20729 11781 20763 11815
rect 3157 11713 3191 11747
rect 4169 11713 4203 11747
rect 10618 11713 10652 11747
rect 10885 11713 10919 11747
rect 11805 11713 11839 11747
rect 20453 11713 20487 11747
rect 1777 11645 1811 11679
rect 1961 11645 1995 11679
rect 2881 11645 2915 11679
rect 4445 11645 4479 11679
rect 5733 11645 5767 11679
rect 5917 11645 5951 11679
rect 7113 11645 7147 11679
rect 7941 11645 7975 11679
rect 14933 11645 14967 11679
rect 17969 11645 18003 11679
rect 3801 11577 3835 11611
rect 19349 11577 19383 11611
rect 6469 11509 6503 11543
rect 7665 11509 7699 11543
rect 9137 11509 9171 11543
rect 16313 11509 16347 11543
rect 16681 11509 16715 11543
rect 20177 11509 20211 11543
rect 3433 11305 3467 11339
rect 9229 11305 9263 11339
rect 10977 11305 11011 11339
rect 11345 11305 11379 11339
rect 15485 11305 15519 11339
rect 19349 11305 19383 11339
rect 21281 11305 21315 11339
rect 5365 11237 5399 11271
rect 13645 11237 13679 11271
rect 2237 11169 2271 11203
rect 2421 11169 2455 11203
rect 3801 11169 3835 11203
rect 4813 11169 4847 11203
rect 6101 11169 6135 11203
rect 6285 11169 6319 11203
rect 7113 11169 7147 11203
rect 7297 11169 7331 11203
rect 8493 11169 8527 11203
rect 10609 11169 10643 11203
rect 2145 11101 2179 11135
rect 7021 11101 7055 11135
rect 8309 11101 8343 11135
rect 10342 11101 10376 11135
rect 14105 11101 14139 11135
rect 14361 11101 14395 11135
rect 16589 11101 16623 11135
rect 18245 11101 18279 11135
rect 18797 11101 18831 11135
rect 20729 11101 20763 11135
rect 1501 11033 1535 11067
rect 4353 11033 4387 11067
rect 4905 11033 4939 11067
rect 6009 11033 6043 11067
rect 8217 11033 8251 11067
rect 16856 11033 16890 11067
rect 20484 11033 20518 11067
rect 1777 10965 1811 10999
rect 2789 10965 2823 10999
rect 4997 10965 5031 10999
rect 5641 10965 5675 10999
rect 6653 10965 6687 10999
rect 7849 10965 7883 10999
rect 15761 10965 15795 10999
rect 17969 10965 18003 10999
rect 1685 10761 1719 10795
rect 2145 10761 2179 10795
rect 2697 10761 2731 10795
rect 3065 10761 3099 10795
rect 3801 10761 3835 10795
rect 4997 10761 5031 10795
rect 6837 10761 6871 10795
rect 7481 10761 7515 10795
rect 9229 10761 9263 10795
rect 15485 10761 15519 10795
rect 19257 10761 19291 10795
rect 21189 10761 21223 10795
rect 2053 10693 2087 10727
rect 18122 10693 18156 10727
rect 19800 10693 19834 10727
rect 5549 10625 5583 10659
rect 7849 10625 7883 10659
rect 10353 10625 10387 10659
rect 14372 10625 14406 10659
rect 17877 10625 17911 10659
rect 2237 10557 2271 10591
rect 3157 10557 3191 10591
rect 3249 10557 3283 10591
rect 6653 10557 6687 10591
rect 6745 10557 6779 10591
rect 7941 10557 7975 10591
rect 8125 10557 8159 10591
rect 8493 10557 8527 10591
rect 10609 10557 10643 10591
rect 10885 10557 10919 10591
rect 11529 10557 11563 10591
rect 14105 10557 14139 10591
rect 19533 10557 19567 10591
rect 5365 10489 5399 10523
rect 20913 10489 20947 10523
rect 4353 10421 4387 10455
rect 5917 10421 5951 10455
rect 7205 10421 7239 10455
rect 8953 10421 8987 10455
rect 15761 10421 15795 10455
rect 1593 10217 1627 10251
rect 7297 10217 7331 10251
rect 10701 10217 10735 10251
rect 16589 10217 16623 10251
rect 20453 10217 20487 10251
rect 2881 10081 2915 10115
rect 5089 10081 5123 10115
rect 5733 10081 5767 10115
rect 7941 10081 7975 10115
rect 21005 10081 21039 10115
rect 3433 10013 3467 10047
rect 4813 10013 4847 10047
rect 6653 10013 6687 10047
rect 9045 10013 9079 10047
rect 12081 10013 12115 10047
rect 14105 10013 14139 10047
rect 15485 10013 15519 10047
rect 18613 10013 18647 10047
rect 19257 10013 19291 10047
rect 19625 10013 19659 10047
rect 2053 9945 2087 9979
rect 2697 9945 2731 9979
rect 7021 9945 7055 9979
rect 9312 9945 9346 9979
rect 11814 9945 11848 9979
rect 16957 9945 16991 9979
rect 18346 9945 18380 9979
rect 2329 9877 2363 9911
rect 2789 9877 2823 9911
rect 4169 9877 4203 9911
rect 4445 9877 4479 9911
rect 4905 9877 4939 9911
rect 6193 9877 6227 9911
rect 7665 9877 7699 9911
rect 7757 9877 7791 9911
rect 8401 9877 8435 9911
rect 10425 9877 10459 9911
rect 12449 9877 12483 9911
rect 17233 9877 17267 9911
rect 20085 9877 20119 9911
rect 20821 9877 20855 9911
rect 20913 9877 20947 9911
rect 5457 9673 5491 9707
rect 11161 9673 11195 9707
rect 14013 9673 14047 9707
rect 21189 9673 21223 9707
rect 1409 9605 1443 9639
rect 7389 9605 7423 9639
rect 9260 9605 9294 9639
rect 10048 9605 10082 9639
rect 12602 9605 12636 9639
rect 16948 9605 16982 9639
rect 19472 9605 19506 9639
rect 20729 9605 20763 9639
rect 3249 9537 3283 9571
rect 4445 9537 4479 9571
rect 5549 9537 5583 9571
rect 7297 9537 7331 9571
rect 15126 9537 15160 9571
rect 15669 9537 15703 9571
rect 20821 9537 20855 9571
rect 2973 9469 3007 9503
rect 3157 9469 3191 9503
rect 4261 9469 4295 9503
rect 4353 9469 4387 9503
rect 5273 9469 5307 9503
rect 7573 9469 7607 9503
rect 9505 9469 9539 9503
rect 9781 9469 9815 9503
rect 12357 9469 12391 9503
rect 15393 9469 15427 9503
rect 15945 9469 15979 9503
rect 16681 9469 16715 9503
rect 19717 9469 19751 9503
rect 19993 9469 20027 9503
rect 20545 9469 20579 9503
rect 1869 9401 1903 9435
rect 3617 9401 3651 9435
rect 4813 9401 4847 9435
rect 8125 9401 8159 9435
rect 11621 9401 11655 9435
rect 18061 9401 18095 9435
rect 2145 9333 2179 9367
rect 2605 9333 2639 9367
rect 5917 9333 5951 9367
rect 6561 9333 6595 9367
rect 6929 9333 6963 9367
rect 13737 9333 13771 9367
rect 18337 9333 18371 9367
rect 1501 9129 1535 9163
rect 3341 9129 3375 9163
rect 10793 9129 10827 9163
rect 13553 9129 13587 9163
rect 14105 9129 14139 9163
rect 3893 8993 3927 9027
rect 4353 8993 4387 9027
rect 5457 8993 5491 9027
rect 5549 8993 5583 9027
rect 6837 8993 6871 9027
rect 8125 8993 8159 9027
rect 11805 8993 11839 9027
rect 18797 8993 18831 9027
rect 19901 8993 19935 9027
rect 20821 8993 20855 9027
rect 20913 8993 20947 9027
rect 2789 8925 2823 8959
rect 4629 8925 4663 8959
rect 6653 8925 6687 8959
rect 7941 8925 7975 8959
rect 9413 8925 9447 8959
rect 11069 8925 11103 8959
rect 12173 8925 12207 8959
rect 12429 8925 12463 8959
rect 15218 8925 15252 8959
rect 15485 8925 15519 8959
rect 15761 8925 15795 8959
rect 16028 8925 16062 8959
rect 19809 8925 19843 8959
rect 2421 8857 2455 8891
rect 5641 8857 5675 8891
rect 6745 8857 6779 8891
rect 9658 8857 9692 8891
rect 17509 8857 17543 8891
rect 18153 8857 18187 8891
rect 19717 8857 19751 8891
rect 4537 8789 4571 8823
rect 4997 8789 5031 8823
rect 6009 8789 6043 8823
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 8033 8789 8067 8823
rect 9045 8789 9079 8823
rect 17141 8789 17175 8823
rect 17785 8789 17819 8823
rect 19349 8789 19383 8823
rect 20361 8789 20395 8823
rect 20729 8789 20763 8823
rect 1869 8585 1903 8619
rect 2329 8585 2363 8619
rect 4537 8585 4571 8619
rect 5549 8585 5583 8619
rect 8033 8585 8067 8619
rect 8125 8585 8159 8619
rect 16773 8585 16807 8619
rect 17877 8585 17911 8619
rect 4997 8517 5031 8551
rect 7021 8517 7055 8551
rect 9137 8517 9171 8551
rect 19266 8517 19300 8551
rect 1961 8449 1995 8483
rect 4261 8449 4295 8483
rect 4905 8449 4939 8483
rect 15229 8449 15263 8483
rect 19533 8449 19567 8483
rect 20922 8449 20956 8483
rect 21189 8449 21223 8483
rect 1777 8381 1811 8415
rect 2789 8381 2823 8415
rect 3801 8381 3835 8415
rect 5181 8381 5215 8415
rect 7941 8381 7975 8415
rect 15485 8381 15519 8415
rect 3249 8313 3283 8347
rect 6561 8313 6595 8347
rect 14105 8313 14139 8347
rect 19809 8313 19843 8347
rect 8493 8245 8527 8279
rect 8769 8245 8803 8279
rect 9689 8245 9723 8279
rect 10425 8245 10459 8279
rect 13645 8245 13679 8279
rect 15853 8245 15887 8279
rect 16129 8245 16163 8279
rect 18153 8245 18187 8279
rect 2237 8041 2271 8075
rect 4169 8041 4203 8075
rect 7665 8041 7699 8075
rect 8953 8041 8987 8075
rect 17969 8041 18003 8075
rect 18797 8041 18831 8075
rect 19993 8041 20027 8075
rect 21005 8041 21039 8075
rect 3801 7973 3835 8007
rect 17233 7973 17267 8007
rect 21281 7973 21315 8007
rect 1685 7905 1719 7939
rect 1777 7905 1811 7939
rect 2697 7905 2731 7939
rect 5549 7905 5583 7939
rect 5733 7905 5767 7939
rect 7113 7905 7147 7939
rect 7297 7905 7331 7939
rect 8217 7905 8251 7939
rect 15853 7905 15887 7939
rect 19349 7905 19383 7939
rect 20361 7905 20395 7939
rect 20545 7905 20579 7939
rect 2881 7837 2915 7871
rect 4905 7837 4939 7871
rect 10066 7837 10100 7871
rect 10333 7837 10367 7871
rect 11722 7837 11756 7871
rect 11989 7837 12023 7871
rect 16109 7837 16143 7871
rect 19533 7837 19567 7871
rect 2789 7769 2823 7803
rect 8033 7769 8067 7803
rect 19625 7769 19659 7803
rect 1869 7701 1903 7735
rect 3249 7701 3283 7735
rect 5825 7701 5859 7735
rect 6193 7701 6227 7735
rect 6653 7701 6687 7735
rect 7021 7701 7055 7735
rect 8125 7701 8159 7735
rect 10609 7701 10643 7735
rect 12265 7701 12299 7735
rect 17509 7701 17543 7735
rect 18521 7701 18555 7735
rect 20637 7701 20671 7735
rect 1593 7497 1627 7531
rect 2329 7497 2363 7531
rect 3341 7497 3375 7531
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 4445 7497 4479 7531
rect 6009 7497 6043 7531
rect 8953 7497 8987 7531
rect 16681 7497 16715 7531
rect 19441 7497 19475 7531
rect 20177 7497 20211 7531
rect 21281 7497 21315 7531
rect 5641 7429 5675 7463
rect 3433 7361 3467 7395
rect 7941 7361 7975 7395
rect 10526 7361 10560 7395
rect 12653 7361 12687 7395
rect 13912 7361 13946 7395
rect 17805 7361 17839 7395
rect 18061 7361 18095 7395
rect 18337 7361 18371 7395
rect 19533 7361 19567 7395
rect 20545 7361 20579 7395
rect 20637 7361 20671 7395
rect 2053 7293 2087 7327
rect 2237 7293 2271 7327
rect 3617 7293 3651 7327
rect 4629 7293 4663 7327
rect 5365 7293 5399 7327
rect 5549 7293 5583 7327
rect 8217 7293 8251 7327
rect 10793 7293 10827 7327
rect 12909 7293 12943 7327
rect 13645 7293 13679 7327
rect 18705 7293 18739 7327
rect 19349 7293 19383 7327
rect 20729 7293 20763 7327
rect 15301 7225 15335 7259
rect 15761 7225 15795 7259
rect 19901 7225 19935 7259
rect 2697 7157 2731 7191
rect 2973 7157 3007 7191
rect 6929 7157 6963 7191
rect 7297 7157 7331 7191
rect 7665 7157 7699 7191
rect 9413 7157 9447 7191
rect 11069 7157 11103 7191
rect 11529 7157 11563 7191
rect 13277 7157 13311 7191
rect 15025 7157 15059 7191
rect 16221 7157 16255 7191
rect 2421 6953 2455 6987
rect 7481 6953 7515 6987
rect 9229 6953 9263 6987
rect 12081 6885 12115 6919
rect 3065 6817 3099 6851
rect 4813 6817 4847 6851
rect 5641 6817 5675 6851
rect 5825 6817 5859 6851
rect 6653 6817 6687 6851
rect 7941 6817 7975 6851
rect 8033 6817 8067 6851
rect 17601 6817 17635 6851
rect 21189 6817 21223 6851
rect 1501 6749 1535 6783
rect 4629 6749 4663 6783
rect 6745 6749 6779 6783
rect 10342 6749 10376 6783
rect 10609 6749 10643 6783
rect 13461 6749 13495 6783
rect 14105 6749 14139 6783
rect 14565 6749 14599 6783
rect 16221 6749 16255 6783
rect 17325 6749 17359 6783
rect 17417 6749 17451 6783
rect 19993 6749 20027 6783
rect 2789 6681 2823 6715
rect 5549 6681 5583 6715
rect 8585 6681 8619 6715
rect 13194 6681 13228 6715
rect 14832 6681 14866 6715
rect 16681 6681 16715 6715
rect 18797 6681 18831 6715
rect 20361 6681 20395 6715
rect 21005 6681 21039 6715
rect 2145 6613 2179 6647
rect 2881 6613 2915 6647
rect 3801 6613 3835 6647
rect 4169 6613 4203 6647
rect 4537 6613 4571 6647
rect 5181 6613 5215 6647
rect 6837 6613 6871 6647
rect 7205 6613 7239 6647
rect 7849 6613 7883 6647
rect 10977 6613 11011 6647
rect 15945 6613 15979 6647
rect 16957 6613 16991 6647
rect 18153 6613 18187 6647
rect 18429 6613 18463 6647
rect 19349 6613 19383 6647
rect 20637 6613 20671 6647
rect 21097 6613 21131 6647
rect 1593 6409 1627 6443
rect 2605 6409 2639 6443
rect 3065 6409 3099 6443
rect 4905 6409 4939 6443
rect 5733 6409 5767 6443
rect 7941 6409 7975 6443
rect 13461 6409 13495 6443
rect 16313 6409 16347 6443
rect 17417 6409 17451 6443
rect 18981 6409 19015 6443
rect 8493 6341 8527 6375
rect 15945 6341 15979 6375
rect 18705 6341 18739 6375
rect 1961 6273 1995 6307
rect 2973 6273 3007 6307
rect 4261 6273 4295 6307
rect 5641 6273 5675 6307
rect 6929 6273 6963 6307
rect 7573 6273 7607 6307
rect 8585 6273 8619 6307
rect 12337 6273 12371 6307
rect 14565 6273 14599 6307
rect 17049 6273 17083 6307
rect 20094 6273 20128 6307
rect 20361 6273 20395 6307
rect 21005 6273 21039 6307
rect 21097 6273 21131 6307
rect 2053 6205 2087 6239
rect 2237 6205 2271 6239
rect 3249 6205 3283 6239
rect 5917 6205 5951 6239
rect 7389 6205 7423 6239
rect 7481 6205 7515 6239
rect 8401 6205 8435 6239
rect 12081 6205 12115 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 16773 6205 16807 6239
rect 16957 6205 16991 6239
rect 21189 6205 21223 6239
rect 8953 6137 8987 6171
rect 14933 6137 14967 6171
rect 3801 6069 3835 6103
rect 4629 6069 4663 6103
rect 5273 6069 5307 6103
rect 6469 6069 6503 6103
rect 9229 6069 9263 6103
rect 9597 6069 9631 6103
rect 13737 6069 13771 6103
rect 15301 6069 15335 6103
rect 17969 6069 18003 6103
rect 18337 6069 18371 6103
rect 20637 6069 20671 6103
rect 4445 5865 4479 5899
rect 5181 5865 5215 5899
rect 5825 5865 5859 5899
rect 21281 5865 21315 5899
rect 5457 5797 5491 5831
rect 9597 5797 9631 5831
rect 21005 5797 21039 5831
rect 1777 5729 1811 5763
rect 3157 5729 3191 5763
rect 3341 5729 3375 5763
rect 6285 5729 6319 5763
rect 6469 5729 6503 5763
rect 8953 5729 8987 5763
rect 13645 5729 13679 5763
rect 18429 5729 18463 5763
rect 19257 5729 19291 5763
rect 4813 5661 4847 5695
rect 6193 5661 6227 5695
rect 8125 5661 8159 5695
rect 10977 5661 11011 5695
rect 15577 5661 15611 5695
rect 17509 5661 17543 5695
rect 17785 5661 17819 5695
rect 2053 5593 2087 5627
rect 3801 5593 3835 5627
rect 7481 5593 7515 5627
rect 8401 5593 8435 5627
rect 10710 5593 10744 5627
rect 15310 5593 15344 5627
rect 17242 5593 17276 5627
rect 19502 5593 19536 5627
rect 1961 5525 1995 5559
rect 2421 5525 2455 5559
rect 2697 5525 2731 5559
rect 3065 5525 3099 5559
rect 7757 5525 7791 5559
rect 11345 5525 11379 5559
rect 11713 5525 11747 5559
rect 14197 5525 14231 5559
rect 16129 5525 16163 5559
rect 18889 5525 18923 5559
rect 20637 5525 20671 5559
rect 2605 5321 2639 5355
rect 3249 5321 3283 5355
rect 4261 5321 4295 5355
rect 4353 5321 4387 5355
rect 8861 5321 8895 5355
rect 15669 5321 15703 5355
rect 16957 5321 16991 5355
rect 17693 5321 17727 5355
rect 20269 5321 20303 5355
rect 21005 5321 21039 5355
rect 5457 5253 5491 5287
rect 13584 5253 13618 5287
rect 15393 5253 15427 5287
rect 20913 5253 20947 5287
rect 5365 5185 5399 5219
rect 6377 5185 6411 5219
rect 7113 5185 7147 5219
rect 8125 5185 8159 5219
rect 9413 5185 9447 5219
rect 9680 5185 9714 5219
rect 11069 5185 11103 5219
rect 13829 5185 13863 5219
rect 14105 5185 14139 5219
rect 14933 5185 14967 5219
rect 17325 5185 17359 5219
rect 18521 5185 18555 5219
rect 19901 5185 19935 5219
rect 1593 5117 1627 5151
rect 2421 5117 2455 5151
rect 2513 5117 2547 5151
rect 4169 5117 4203 5151
rect 5641 5117 5675 5151
rect 7389 5117 7423 5151
rect 8309 5117 8343 5151
rect 19625 5117 19659 5151
rect 19809 5117 19843 5151
rect 21097 5117 21131 5151
rect 12449 5049 12483 5083
rect 16221 5049 16255 5083
rect 18153 5049 18187 5083
rect 18889 5049 18923 5083
rect 20545 5049 20579 5083
rect 1869 4981 1903 5015
rect 2973 4981 3007 5015
rect 3709 4981 3743 5015
rect 4721 4981 4755 5015
rect 4997 4981 5031 5015
rect 10793 4981 10827 5015
rect 11805 4981 11839 5015
rect 14657 4981 14691 5015
rect 19165 4981 19199 5015
rect 1777 4777 1811 4811
rect 2145 4777 2179 4811
rect 3249 4777 3283 4811
rect 6377 4777 6411 4811
rect 9689 4777 9723 4811
rect 12265 4777 12299 4811
rect 15485 4777 15519 4811
rect 17141 4777 17175 4811
rect 20637 4777 20671 4811
rect 20913 4777 20947 4811
rect 10333 4709 10367 4743
rect 2697 4641 2731 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 5825 4641 5859 4675
rect 5917 4641 5951 4675
rect 9137 4641 9171 4675
rect 9229 4641 9263 4675
rect 10057 4641 10091 4675
rect 13645 4641 13679 4675
rect 14105 4641 14139 4675
rect 19257 4641 19291 4675
rect 1501 4573 1535 4607
rect 2881 4573 2915 4607
rect 4261 4573 4295 4607
rect 4905 4573 4939 4607
rect 6653 4573 6687 4607
rect 8033 4573 8067 4607
rect 11713 4573 11747 4607
rect 16609 4573 16643 4607
rect 16865 4573 16899 4607
rect 18521 4573 18555 4607
rect 18797 4573 18831 4607
rect 6009 4505 6043 4539
rect 6929 4505 6963 4539
rect 8309 4505 8343 4539
rect 11446 4505 11480 4539
rect 13378 4505 13412 4539
rect 14841 4505 14875 4539
rect 18276 4505 18310 4539
rect 19524 4505 19558 4539
rect 2789 4437 2823 4471
rect 3893 4437 3927 4471
rect 5273 4437 5307 4471
rect 7757 4437 7791 4471
rect 9321 4437 9355 4471
rect 15209 4437 15243 4471
rect 21373 4437 21407 4471
rect 3801 4233 3835 4267
rect 7941 4233 7975 4267
rect 8953 4233 8987 4267
rect 17509 4233 17543 4267
rect 18613 4233 18647 4267
rect 3893 4165 3927 4199
rect 10894 4165 10928 4199
rect 16221 4165 16255 4199
rect 2513 4097 2547 4131
rect 3157 4097 3191 4131
rect 6377 4097 6411 4131
rect 7481 4097 7515 4131
rect 8861 4097 8895 4131
rect 11161 4097 11195 4131
rect 11529 4097 11563 4131
rect 13093 4097 13127 4131
rect 13461 4097 13495 4131
rect 15310 4097 15344 4131
rect 15577 4097 15611 4131
rect 20462 4097 20496 4131
rect 20729 4097 20763 4131
rect 21281 4097 21315 4131
rect 2329 4029 2363 4063
rect 2421 4029 2455 4063
rect 3709 4029 3743 4063
rect 6653 4029 6687 4063
rect 8769 4029 8803 4063
rect 17601 4029 17635 4063
rect 17693 4029 17727 4063
rect 18981 4029 19015 4063
rect 8309 3961 8343 3995
rect 9321 3961 9355 3995
rect 9781 3961 9815 3995
rect 11989 3961 12023 3995
rect 15945 3961 15979 3995
rect 17141 3961 17175 3995
rect 18153 3961 18187 3995
rect 1409 3893 1443 3927
rect 1777 3893 1811 3927
rect 2881 3893 2915 3927
rect 4261 3893 4295 3927
rect 5917 3893 5951 3927
rect 7205 3893 7239 3927
rect 12357 3893 12391 3927
rect 13737 3893 13771 3927
rect 14197 3893 14231 3927
rect 16865 3893 16899 3927
rect 19349 3893 19383 3927
rect 21097 3893 21131 3927
rect 2605 3689 2639 3723
rect 3433 3689 3467 3723
rect 8125 3689 8159 3723
rect 10609 3689 10643 3723
rect 12265 3689 12299 3723
rect 14381 3689 14415 3723
rect 16313 3689 16347 3723
rect 17877 3689 17911 3723
rect 20361 3689 20395 3723
rect 1593 3621 1627 3655
rect 6745 3621 6779 3655
rect 7205 3621 7239 3655
rect 15945 3621 15979 3655
rect 16773 3621 16807 3655
rect 19901 3621 19935 3655
rect 1961 3553 1995 3587
rect 2145 3553 2179 3587
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 6193 3553 6227 3587
rect 9597 3553 9631 3587
rect 11982 3553 12016 3587
rect 15025 3553 15059 3587
rect 15485 3553 15519 3587
rect 17325 3553 17359 3587
rect 17417 3553 17451 3587
rect 18797 3553 18831 3587
rect 19257 3553 19291 3587
rect 20913 3553 20947 3587
rect 4261 3485 4295 3519
rect 4997 3485 5031 3519
rect 7021 3485 7055 3519
rect 7573 3485 7607 3519
rect 13645 3485 13679 3519
rect 16589 3485 16623 3519
rect 18613 3485 18647 3519
rect 20085 3485 20119 3519
rect 20729 3485 20763 3519
rect 20821 3485 20855 3519
rect 6285 3417 6319 3451
rect 10333 3417 10367 3451
rect 11744 3417 11778 3451
rect 13378 3417 13412 3451
rect 14749 3417 14783 3451
rect 14841 3417 14875 3451
rect 18521 3417 18555 3451
rect 2237 3349 2271 3383
rect 2881 3349 2915 3383
rect 3893 3349 3927 3383
rect 5733 3349 5767 3383
rect 6377 3349 6411 3383
rect 7757 3349 7791 3383
rect 8585 3349 8619 3383
rect 8953 3349 8987 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 17509 3349 17543 3383
rect 18153 3349 18187 3383
rect 4353 3145 4387 3179
rect 4813 3145 4847 3179
rect 6837 3145 6871 3179
rect 7849 3145 7883 3179
rect 12633 3145 12667 3179
rect 13277 3145 13311 3179
rect 13645 3145 13679 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 17693 3145 17727 3179
rect 18061 3145 18095 3179
rect 19073 3145 19107 3179
rect 21373 3145 21407 3179
rect 2973 3077 3007 3111
rect 4721 3077 4755 3111
rect 5641 3077 5675 3111
rect 6745 3077 6779 3111
rect 11529 3077 11563 3111
rect 12173 3077 12207 3111
rect 14197 3077 14231 3111
rect 16129 3077 16163 3111
rect 19165 3077 19199 3111
rect 20821 3077 20855 3111
rect 1961 3009 1995 3043
rect 2513 3009 2547 3043
rect 3801 3009 3835 3043
rect 4077 3009 4111 3043
rect 7665 3009 7699 3043
rect 8217 3009 8251 3043
rect 9229 3009 9263 3043
rect 10894 3009 10928 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 13921 3009 13955 3043
rect 14841 3009 14875 3043
rect 15577 3009 15611 3043
rect 18153 3009 18187 3043
rect 19993 3009 20027 3043
rect 4997 2941 5031 2975
rect 7021 2941 7055 2975
rect 9045 2941 9079 2975
rect 12081 2941 12115 2975
rect 13001 2941 13035 2975
rect 13185 2941 13219 2975
rect 15117 2941 15151 2975
rect 17141 2941 17175 2975
rect 17233 2941 17267 2975
rect 18337 2941 18371 2975
rect 19257 2941 19291 2975
rect 6377 2873 6411 2907
rect 8401 2873 8435 2907
rect 15761 2873 15795 2907
rect 18705 2873 18739 2907
rect 2145 2805 2179 2839
rect 3249 2805 3283 2839
rect 6009 2805 6043 2839
rect 9781 2805 9815 2839
rect 4077 2601 4111 2635
rect 5181 2601 5215 2635
rect 9781 2601 9815 2635
rect 12541 2601 12575 2635
rect 12909 2601 12943 2635
rect 14197 2601 14231 2635
rect 14565 2601 14599 2635
rect 18521 2601 18555 2635
rect 20637 2601 20671 2635
rect 19349 2533 19383 2567
rect 4629 2465 4663 2499
rect 5641 2465 5675 2499
rect 6745 2465 6779 2499
rect 13369 2465 13403 2499
rect 13553 2465 13587 2499
rect 16957 2465 16991 2499
rect 21189 2465 21223 2499
rect 5917 2397 5951 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7849 2397 7883 2431
rect 8953 2397 8987 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 11713 2397 11747 2431
rect 15117 2397 15151 2431
rect 15761 2397 15795 2431
rect 17141 2397 17175 2431
rect 17417 2397 17451 2431
rect 18245 2397 18279 2431
rect 19533 2397 19567 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 4537 2329 4571 2363
rect 13277 2329 13311 2363
rect 3433 2261 3467 2295
rect 4445 2261 4479 2295
rect 7389 2261 7423 2295
rect 8033 2261 8067 2295
rect 8585 2261 8619 2295
rect 9137 2261 9171 2295
rect 10241 2261 10275 2295
rect 10885 2261 10919 2295
rect 11897 2261 11931 2295
rect 15301 2261 15335 2295
rect 15945 2261 15979 2295
rect 17601 2261 17635 2295
rect 18061 2261 18095 2295
rect 20269 2261 20303 2295
rect 21097 2261 21131 2295
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20312 20556 21005 20584
rect 20312 20544 20318 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 13722 20476 13728 20528
rect 13780 20516 13786 20528
rect 13780 20488 17172 20516
rect 13780 20476 13786 20488
rect 2133 20451 2191 20457
rect 2133 20417 2145 20451
rect 2179 20448 2191 20451
rect 14093 20451 14151 20457
rect 2179 20420 2544 20448
rect 2179 20417 2191 20420
rect 2133 20411 2191 20417
rect 2516 20253 2544 20420
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14366 20448 14372 20460
rect 14139 20420 14372 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 7834 20380 7840 20392
rect 7795 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 17144 20389 17172 20488
rect 17773 20451 17831 20457
rect 17773 20417 17785 20451
rect 17819 20448 17831 20451
rect 18230 20448 18236 20460
rect 17819 20420 18236 20448
rect 17819 20417 17831 20420
rect 17773 20411 17831 20417
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 19886 20408 19892 20460
rect 19944 20448 19950 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 19944 20420 20269 20448
rect 19944 20408 19950 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17175 20352 17877 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 17865 20349 17877 20352
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 18138 20380 18144 20392
rect 18095 20352 18144 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 14292 20312 14320 20343
rect 18138 20340 18144 20352
rect 18196 20340 18202 20392
rect 20824 20312 20852 20411
rect 14292 20284 20852 20312
rect 2501 20247 2559 20253
rect 2501 20213 2513 20247
rect 2547 20244 2559 20247
rect 4062 20244 4068 20256
rect 2547 20216 4068 20244
rect 2547 20213 2559 20216
rect 2501 20207 2559 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 12342 20244 12348 20256
rect 12303 20216 12348 20244
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 17402 20244 17408 20256
rect 17363 20216 17408 20244
rect 17402 20204 17408 20216
rect 17460 20204 17466 20256
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 18417 20247 18475 20253
rect 18417 20244 18429 20247
rect 18196 20216 18429 20244
rect 18196 20204 18202 20216
rect 18417 20213 18429 20216
rect 18463 20213 18475 20247
rect 18417 20207 18475 20213
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 19886 20244 19892 20256
rect 18564 20216 19892 20244
rect 18564 20204 18570 20216
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 20438 20244 20444 20256
rect 20399 20216 20444 20244
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 2774 20040 2780 20052
rect 2547 20012 2780 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 13722 20040 13728 20052
rect 13683 20012 13728 20040
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14093 20043 14151 20049
rect 14093 20009 14105 20043
rect 14139 20040 14151 20043
rect 14366 20040 14372 20052
rect 14139 20012 14372 20040
rect 14139 20009 14151 20012
rect 14093 20003 14151 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 18046 20040 18052 20052
rect 14608 20012 18052 20040
rect 14608 20000 14614 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 20680 20012 20913 20040
rect 20680 20000 20686 20012
rect 20901 20009 20913 20012
rect 20947 20009 20959 20043
rect 20901 20003 20959 20009
rect 12618 19972 12624 19984
rect 11992 19944 12624 19972
rect 3973 19907 4031 19913
rect 3973 19904 3985 19907
rect 2148 19876 3985 19904
rect 2148 19845 2176 19876
rect 3973 19873 3985 19876
rect 4019 19873 4031 19907
rect 3973 19867 4031 19873
rect 7653 19907 7711 19913
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 8478 19904 8484 19916
rect 7699 19876 8484 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 10502 19904 10508 19916
rect 10463 19876 10508 19904
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 10888 19876 11897 19904
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2731 19808 2973 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 2961 19805 2973 19808
rect 3007 19836 3019 19839
rect 3878 19836 3884 19848
rect 3007 19808 3884 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 4706 19836 4712 19848
rect 4295 19808 4712 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 10888 19836 10916 19876
rect 11885 19873 11897 19876
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 9916 19808 10916 19836
rect 9916 19796 9922 19808
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11112 19808 11805 19836
rect 11112 19796 11118 19808
rect 11793 19805 11805 19808
rect 11839 19836 11851 19839
rect 11992 19836 12020 19944
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 12713 19975 12771 19981
rect 12713 19941 12725 19975
rect 12759 19972 12771 19975
rect 17954 19972 17960 19984
rect 12759 19944 17960 19972
rect 12759 19941 12771 19944
rect 12713 19935 12771 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 13722 19904 13728 19916
rect 12492 19876 13728 19904
rect 12492 19864 12498 19876
rect 11839 19808 12020 19836
rect 11839 19805 11851 19808
rect 11793 19799 11851 19805
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 13096 19845 13124 19876
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 14734 19904 14740 19916
rect 14695 19876 14740 19904
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16080 19876 16681 19904
rect 16080 19864 16086 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19904 17371 19907
rect 17678 19904 17684 19916
rect 17359 19876 17684 19904
rect 17359 19873 17371 19876
rect 17313 19867 17371 19873
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 18230 19904 18236 19916
rect 18191 19876 18236 19904
rect 18230 19864 18236 19876
rect 18288 19864 18294 19916
rect 12529 19839 12587 19845
rect 12529 19836 12541 19839
rect 12400 19808 12541 19836
rect 12400 19796 12434 19808
rect 12529 19805 12541 19808
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13630 19796 13636 19848
rect 13688 19836 13694 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 13688 19808 14565 19836
rect 13688 19796 13694 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 14884 19808 15117 19836
rect 14884 19796 14890 19808
rect 15105 19805 15117 19808
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 17402 19836 17408 19848
rect 16531 19808 17408 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 17972 19808 19257 19836
rect 10321 19771 10379 19777
rect 10321 19737 10333 19771
rect 10367 19768 10379 19771
rect 10367 19740 11376 19768
rect 10367 19737 10379 19740
rect 10321 19731 10379 19737
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 7098 19700 7104 19712
rect 7059 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19700 7162 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7156 19672 7757 19700
rect 7156 19660 7162 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7984 19672 8217 19700
rect 7984 19660 7990 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 9950 19700 9956 19712
rect 9911 19672 9956 19700
rect 8205 19663 8263 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 11054 19700 11060 19712
rect 10468 19672 10513 19700
rect 11015 19672 11060 19700
rect 10468 19660 10474 19672
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11348 19709 11376 19740
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 12406 19768 12434 19796
rect 11940 19740 12434 19768
rect 14461 19771 14519 19777
rect 11940 19728 11946 19740
rect 14461 19737 14473 19771
rect 14507 19768 14519 19771
rect 14507 19740 15148 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 11333 19703 11391 19709
rect 11333 19669 11345 19703
rect 11379 19669 11391 19703
rect 11698 19700 11704 19712
rect 11659 19672 11704 19700
rect 11333 19663 11391 19669
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 13265 19703 13323 19709
rect 13265 19669 13277 19703
rect 13311 19700 13323 19703
rect 14550 19700 14556 19712
rect 13311 19672 14556 19700
rect 13311 19669 13323 19672
rect 13265 19663 13323 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 15120 19700 15148 19740
rect 15378 19728 15384 19780
rect 15436 19768 15442 19780
rect 15436 19740 15481 19768
rect 15436 19728 15442 19740
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15120 19672 16129 19700
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16942 19700 16948 19712
rect 16623 19672 16948 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17494 19700 17500 19712
rect 17455 19672 17500 19700
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 17972 19709 18000 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19567 19808 19993 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 20714 19836 20720 19848
rect 20675 19808 20720 19836
rect 19981 19799 20039 19805
rect 20714 19796 20720 19808
rect 20772 19836 20778 19848
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 20772 19808 21281 19836
rect 20772 19796 20778 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 17957 19703 18015 19709
rect 17644 19672 17689 19700
rect 17644 19660 17650 19672
rect 17957 19669 17969 19703
rect 18003 19669 18015 19703
rect 18690 19700 18696 19712
rect 18651 19672 18696 19700
rect 17957 19663 18015 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2501 19499 2559 19505
rect 2501 19465 2513 19499
rect 2547 19496 2559 19499
rect 2866 19496 2872 19508
rect 2547 19468 2872 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 7926 19496 7932 19508
rect 7887 19468 7932 19496
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 10410 19496 10416 19508
rect 10371 19468 10416 19496
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11756 19468 11805 19496
rect 11756 19456 11762 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 12618 19456 12624 19508
rect 12676 19496 12682 19508
rect 14826 19496 14832 19508
rect 12676 19468 14688 19496
rect 14787 19468 14832 19496
rect 12676 19456 12682 19468
rect 14366 19428 14372 19440
rect 14327 19400 14372 19428
rect 14366 19388 14372 19400
rect 14424 19388 14430 19440
rect 14660 19428 14688 19468
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 16022 19496 16028 19508
rect 15983 19468 16028 19496
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 17126 19496 17132 19508
rect 17087 19468 17132 19496
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17586 19496 17592 19508
rect 17451 19468 17592 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 17773 19499 17831 19505
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 18690 19496 18696 19508
rect 17819 19468 18696 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 18506 19428 18512 19440
rect 14660 19400 18512 19428
rect 18506 19388 18512 19400
rect 18564 19388 18570 19440
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1627 19332 2145 19360
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 2133 19329 2145 19332
rect 2179 19360 2191 19363
rect 2498 19360 2504 19372
rect 2179 19332 2504 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 2498 19320 2504 19332
rect 2556 19320 2562 19372
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 5074 19360 5080 19372
rect 2731 19332 3004 19360
rect 5035 19332 5080 19360
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2976 19301 3004 19332
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 5166 19320 5172 19372
rect 5224 19360 5230 19372
rect 5224 19332 5269 19360
rect 5224 19320 5230 19332
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 8628 19332 10057 19360
rect 8628 19320 8634 19332
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3970 19292 3976 19304
rect 3007 19264 3976 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 6457 19295 6515 19301
rect 6457 19261 6469 19295
rect 6503 19292 6515 19295
rect 7282 19292 7288 19304
rect 6503 19264 7288 19292
rect 6503 19261 6515 19264
rect 6457 19255 6515 19261
rect 1946 19224 1952 19236
rect 1907 19196 1952 19224
rect 1946 19184 1952 19196
rect 2004 19184 2010 19236
rect 5368 19224 5396 19255
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 8018 19292 8024 19304
rect 7979 19264 8024 19292
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19292 8263 19295
rect 9306 19292 9312 19304
rect 8251 19264 9312 19292
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 9416 19301 9444 19332
rect 10045 19329 10057 19332
rect 10091 19329 10103 19363
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 10045 19323 10103 19329
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 15436 19332 20729 19360
rect 15436 19320 15442 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 9401 19295 9459 19301
rect 9401 19261 9413 19295
rect 9447 19261 9459 19295
rect 9858 19292 9864 19304
rect 9819 19264 9864 19292
rect 9401 19255 9459 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 10134 19292 10140 19304
rect 9999 19264 10140 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 10134 19252 10140 19264
rect 10192 19292 10198 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 10192 19264 10701 19292
rect 10192 19252 10198 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 12342 19292 12348 19304
rect 12303 19264 12348 19292
rect 10689 19255 10747 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 15470 19292 15476 19304
rect 14323 19264 15476 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 17770 19292 17776 19304
rect 16684 19264 17776 19292
rect 5813 19227 5871 19233
rect 5813 19224 5825 19227
rect 5368 19196 5825 19224
rect 5813 19193 5825 19196
rect 5859 19224 5871 19227
rect 5859 19196 15967 19224
rect 5859 19193 5871 19196
rect 5813 19187 5871 19193
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 6733 19159 6791 19165
rect 6733 19156 6745 19159
rect 6604 19128 6745 19156
rect 6604 19116 6610 19128
rect 6733 19125 6745 19128
rect 6779 19125 6791 19159
rect 7558 19156 7564 19168
rect 7519 19128 7564 19156
rect 6733 19119 6791 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15252 19128 15393 19156
rect 15252 19116 15258 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15939 19156 15967 19196
rect 16482 19184 16488 19236
rect 16540 19224 16546 19236
rect 16684 19233 16712 19264
rect 17770 19252 17776 19264
rect 17828 19292 17834 19304
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17828 19264 17877 19292
rect 17828 19252 17834 19264
rect 17865 19261 17877 19264
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 17957 19295 18015 19301
rect 17957 19261 17969 19295
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 16669 19227 16727 19233
rect 16669 19224 16681 19227
rect 16540 19196 16681 19224
rect 16540 19184 16546 19196
rect 16669 19193 16681 19196
rect 16715 19193 16727 19227
rect 17972 19224 18000 19255
rect 16669 19187 16727 19193
rect 17880 19196 18000 19224
rect 17880 19168 17908 19196
rect 17218 19156 17224 19168
rect 15939 19128 17224 19156
rect 15381 19119 15439 19125
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 17862 19116 17868 19168
rect 17920 19116 17926 19168
rect 20898 19156 20904 19168
rect 20859 19128 20904 19156
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 5132 18924 5273 18952
rect 5132 18912 5138 18924
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 13538 18952 13544 18964
rect 5261 18915 5319 18921
rect 9324 18924 13544 18952
rect 3789 18887 3847 18893
rect 3789 18853 3801 18887
rect 3835 18853 3847 18887
rect 3789 18847 3847 18853
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 3053 18751 3111 18757
rect 3053 18748 3065 18751
rect 2179 18720 3065 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 3053 18717 3065 18720
rect 3099 18717 3111 18751
rect 3053 18711 3111 18717
rect 3329 18751 3387 18757
rect 3329 18717 3341 18751
rect 3375 18748 3387 18751
rect 3804 18748 3832 18847
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 5074 18816 5080 18828
rect 4479 18788 5080 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18816 5963 18819
rect 6546 18816 6552 18828
rect 5951 18788 6552 18816
rect 5951 18785 5963 18788
rect 5905 18779 5963 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 8938 18816 8944 18828
rect 6880 18788 8944 18816
rect 6880 18776 6886 18788
rect 8938 18776 8944 18788
rect 8996 18816 9002 18828
rect 9324 18816 9352 18924
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 14516 18924 14565 18952
rect 14516 18912 14522 18924
rect 14553 18921 14565 18924
rect 14599 18921 14611 18955
rect 14553 18915 14611 18921
rect 14642 18912 14648 18964
rect 14700 18952 14706 18964
rect 16482 18952 16488 18964
rect 14700 18924 16488 18952
rect 14700 18912 14706 18924
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 16577 18955 16635 18961
rect 16577 18921 16589 18955
rect 16623 18952 16635 18955
rect 16942 18952 16948 18964
rect 16623 18924 16948 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18322 18952 18328 18964
rect 17828 18924 18328 18952
rect 17828 18912 17834 18924
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18506 18952 18512 18964
rect 18467 18924 18512 18952
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 12066 18844 12072 18896
rect 12124 18884 12130 18896
rect 12434 18884 12440 18896
rect 12124 18856 12440 18884
rect 12124 18844 12130 18856
rect 12434 18844 12440 18856
rect 12492 18844 12498 18896
rect 18690 18884 18696 18896
rect 15028 18856 18696 18884
rect 8996 18788 9352 18816
rect 8996 18776 9002 18788
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11020 18788 11989 18816
rect 11020 18776 11026 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 12618 18816 12624 18828
rect 12579 18788 12624 18816
rect 11977 18779 12035 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 15028 18816 15056 18856
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 19981 18887 20039 18893
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 20806 18884 20812 18896
rect 20027 18856 20812 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 14936 18788 15056 18816
rect 15105 18819 15163 18825
rect 3375 18720 3832 18748
rect 4157 18751 4215 18757
rect 3375 18717 3387 18720
rect 3329 18711 3387 18717
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 4246 18748 4252 18760
rect 4203 18720 4252 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 7929 18751 7987 18757
rect 7929 18748 7941 18751
rect 5552 18720 7941 18748
rect 1762 18640 1768 18692
rect 1820 18680 1826 18692
rect 5552 18680 5580 18720
rect 7929 18717 7941 18720
rect 7975 18748 7987 18751
rect 8294 18748 8300 18760
rect 7975 18720 8300 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 8294 18708 8300 18720
rect 8352 18748 8358 18760
rect 11606 18748 11612 18760
rect 8352 18720 11612 18748
rect 8352 18708 8358 18720
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 12342 18748 12348 18760
rect 11839 18720 12348 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 14936 18748 14964 18788
rect 15105 18785 15117 18819
rect 15151 18785 15163 18819
rect 16114 18816 16120 18828
rect 16075 18788 16120 18816
rect 15105 18779 15163 18785
rect 13188 18720 14964 18748
rect 1820 18652 5580 18680
rect 5629 18683 5687 18689
rect 1820 18640 1826 18652
rect 5629 18649 5641 18683
rect 5675 18680 5687 18683
rect 6273 18683 6331 18689
rect 6273 18680 6285 18683
rect 5675 18652 6285 18680
rect 5675 18649 5687 18652
rect 5629 18643 5687 18649
rect 6273 18649 6285 18652
rect 6319 18649 6331 18683
rect 7101 18683 7159 18689
rect 7101 18680 7113 18683
rect 6273 18643 6331 18649
rect 6380 18652 7113 18680
rect 1946 18612 1952 18624
rect 1907 18584 1952 18612
rect 1946 18572 1952 18584
rect 2004 18572 2010 18624
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 3142 18612 3148 18624
rect 2639 18584 3148 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4522 18612 4528 18624
rect 4295 18584 4528 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 6380 18612 6408 18652
rect 7101 18649 7113 18652
rect 7147 18649 7159 18683
rect 7101 18643 7159 18649
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 10318 18680 10324 18692
rect 7340 18652 10324 18680
rect 7340 18640 7346 18652
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 11072 18652 11560 18680
rect 11072 18624 11100 18652
rect 5960 18584 6408 18612
rect 5960 18572 5966 18584
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 6604 18584 6745 18612
rect 6604 18572 6610 18584
rect 6733 18581 6745 18584
rect 6779 18581 6791 18615
rect 6733 18575 6791 18581
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 7561 18615 7619 18621
rect 7561 18612 7573 18615
rect 7248 18584 7573 18612
rect 7248 18572 7254 18584
rect 7561 18581 7573 18584
rect 7607 18581 7619 18615
rect 7561 18575 7619 18581
rect 9493 18615 9551 18621
rect 9493 18581 9505 18615
rect 9539 18612 9551 18615
rect 9674 18612 9680 18624
rect 9539 18584 9680 18612
rect 9539 18581 9551 18584
rect 9493 18575 9551 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 9861 18615 9919 18621
rect 9861 18581 9873 18615
rect 9907 18612 9919 18615
rect 9950 18612 9956 18624
rect 9907 18584 9956 18612
rect 9907 18581 9919 18584
rect 9861 18575 9919 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 11054 18612 11060 18624
rect 11015 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11296 18584 11437 18612
rect 11296 18572 11302 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 11532 18612 11560 18652
rect 11698 18640 11704 18692
rect 11756 18680 11762 18692
rect 12713 18683 12771 18689
rect 12713 18680 12725 18683
rect 11756 18652 12725 18680
rect 11756 18640 11762 18652
rect 12713 18649 12725 18652
rect 12759 18649 12771 18683
rect 12713 18643 12771 18649
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 11532 18584 11897 18612
rect 11425 18575 11483 18581
rect 11885 18581 11897 18584
rect 11931 18612 11943 18615
rect 12066 18612 12072 18624
rect 11931 18584 12072 18612
rect 11931 18581 11943 18584
rect 11885 18575 11943 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12802 18612 12808 18624
rect 12763 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 13188 18621 13216 18720
rect 15010 18708 15016 18760
rect 15068 18748 15074 18760
rect 15120 18748 15148 18779
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 17221 18819 17279 18825
rect 17221 18816 17233 18819
rect 17184 18788 17233 18816
rect 17184 18776 17190 18788
rect 17221 18785 17233 18788
rect 17267 18816 17279 18819
rect 18138 18816 18144 18828
rect 17267 18788 18144 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 19521 18819 19579 18825
rect 19521 18785 19533 18819
rect 19567 18816 19579 18819
rect 20162 18816 20168 18828
rect 19567 18788 20168 18816
rect 19567 18785 19579 18788
rect 19521 18779 19579 18785
rect 15068 18720 15148 18748
rect 15068 18708 15074 18720
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15252 18720 15945 18748
rect 15252 18708 15258 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16264 18720 17049 18748
rect 16264 18708 16270 18720
rect 17037 18717 17049 18720
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 18230 18708 18236 18760
rect 18288 18748 18294 18760
rect 18598 18748 18604 18760
rect 18288 18720 18604 18748
rect 18288 18708 18294 18720
rect 18598 18708 18604 18720
rect 18656 18748 18662 18760
rect 19352 18748 19380 18779
rect 20162 18776 20168 18788
rect 20220 18776 20226 18828
rect 18656 18720 19380 18748
rect 18656 18708 18662 18720
rect 19794 18708 19800 18760
rect 19852 18748 19858 18760
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 19852 18720 20821 18748
rect 19852 18708 19858 18720
rect 20809 18717 20821 18720
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 14921 18683 14979 18689
rect 14921 18649 14933 18683
rect 14967 18680 14979 18683
rect 16390 18680 16396 18692
rect 14967 18652 16396 18680
rect 14967 18649 14979 18652
rect 14921 18643 14979 18649
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 16942 18680 16948 18692
rect 16903 18652 16948 18680
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 18104 18652 18149 18680
rect 18104 18640 18110 18652
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18932 18652 21036 18680
rect 18932 18640 18938 18652
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18581 13231 18615
rect 13173 18575 13231 18581
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 15068 18584 15113 18612
rect 15068 18572 15074 18584
rect 15378 18572 15384 18624
rect 15436 18612 15442 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15436 18584 15577 18612
rect 15436 18572 15442 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16080 18584 16125 18612
rect 16080 18572 16086 18584
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17589 18615 17647 18621
rect 17589 18612 17601 18615
rect 17552 18584 17601 18612
rect 17552 18572 17558 18584
rect 17589 18581 17601 18584
rect 17635 18612 17647 18615
rect 19426 18612 19432 18624
rect 17635 18584 19432 18612
rect 17635 18581 17647 18584
rect 17589 18575 17647 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 19610 18612 19616 18624
rect 19571 18584 19616 18612
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 20346 18612 20352 18624
rect 20307 18584 20352 18612
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 21008 18621 21036 18652
rect 20993 18615 21051 18621
rect 20993 18581 21005 18615
rect 21039 18581 21051 18615
rect 20993 18575 21051 18581
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4249 18411 4307 18417
rect 4249 18408 4261 18411
rect 3651 18380 4261 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4249 18377 4261 18380
rect 4295 18377 4307 18411
rect 4249 18371 4307 18377
rect 5721 18411 5779 18417
rect 5721 18377 5733 18411
rect 5767 18408 5779 18411
rect 7282 18408 7288 18420
rect 5767 18380 7288 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 5736 18340 5764 18371
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 7929 18411 7987 18417
rect 7929 18377 7941 18411
rect 7975 18408 7987 18411
rect 8018 18408 8024 18420
rect 7975 18380 8024 18408
rect 7975 18377 7987 18380
rect 7929 18371 7987 18377
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8294 18408 8300 18420
rect 8255 18380 8300 18408
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 10042 18408 10048 18420
rect 8536 18380 10048 18408
rect 8536 18368 8542 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10137 18411 10195 18417
rect 10137 18377 10149 18411
rect 10183 18377 10195 18411
rect 10137 18371 10195 18377
rect 12345 18411 12403 18417
rect 12345 18377 12357 18411
rect 12391 18408 12403 18411
rect 12802 18408 12808 18420
rect 12391 18380 12808 18408
rect 12391 18377 12403 18380
rect 12345 18371 12403 18377
rect 2148 18312 5764 18340
rect 2148 18281 2176 18312
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 6972 18312 7665 18340
rect 6972 18300 6978 18312
rect 7653 18309 7665 18312
rect 7699 18340 7711 18343
rect 10152 18340 10180 18371
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13814 18408 13820 18420
rect 13775 18380 13820 18408
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 15378 18408 15384 18420
rect 15339 18380 15384 18408
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17972 18380 18061 18408
rect 17402 18340 17408 18352
rect 7699 18312 9674 18340
rect 10152 18312 17408 18340
rect 7699 18309 7711 18312
rect 7653 18303 7711 18309
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 1627 18244 2145 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2133 18241 2145 18244
rect 2179 18241 2191 18275
rect 3234 18272 3240 18284
rect 3195 18244 3240 18272
rect 2133 18235 2191 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4985 18275 5043 18281
rect 4985 18272 4997 18275
rect 4120 18244 4997 18272
rect 4120 18232 4126 18244
rect 4985 18241 4997 18244
rect 5031 18272 5043 18275
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5031 18244 5641 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 5629 18241 5641 18244
rect 5675 18272 5687 18275
rect 5994 18272 6000 18284
rect 5675 18244 6000 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 5994 18232 6000 18244
rect 6052 18232 6058 18284
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8662 18272 8668 18284
rect 8435 18244 8668 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 9309 18275 9367 18281
rect 9309 18272 9321 18275
rect 8996 18244 9321 18272
rect 8996 18232 9002 18244
rect 9309 18241 9321 18244
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18173 3019 18207
rect 3142 18204 3148 18216
rect 3103 18176 3148 18204
rect 2961 18167 3019 18173
rect 1578 18028 1584 18080
rect 1636 18068 1642 18080
rect 1949 18071 2007 18077
rect 1949 18068 1961 18071
rect 1636 18040 1961 18068
rect 1636 18028 1642 18040
rect 1949 18037 1961 18040
rect 1995 18037 2007 18071
rect 2406 18068 2412 18080
rect 2367 18040 2412 18068
rect 1949 18031 2007 18037
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 2976 18068 3004 18167
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18173 4031 18207
rect 4154 18204 4160 18216
rect 4115 18176 4160 18204
rect 3973 18167 4031 18173
rect 3988 18136 4016 18167
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 4798 18204 4804 18216
rect 4264 18176 4804 18204
rect 4264 18136 4292 18176
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 5902 18204 5908 18216
rect 5863 18176 5908 18204
rect 5902 18164 5908 18176
rect 5960 18164 5966 18216
rect 8478 18204 8484 18216
rect 8439 18176 8484 18204
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 9398 18204 9404 18216
rect 9359 18176 9404 18204
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 9646 18204 9674 18312
rect 17402 18300 17408 18312
rect 17460 18300 17466 18352
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 17972 18340 18000 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 18141 18411 18199 18417
rect 18141 18377 18153 18411
rect 18187 18408 18199 18411
rect 18506 18408 18512 18420
rect 18187 18380 18512 18408
rect 18187 18377 18199 18380
rect 18141 18371 18199 18377
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 19150 18340 19156 18352
rect 17552 18312 18000 18340
rect 19111 18312 19156 18340
rect 17552 18300 17558 18312
rect 19150 18300 19156 18312
rect 19208 18300 19214 18352
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 19484 18312 20852 18340
rect 19484 18300 19490 18312
rect 9950 18272 9956 18284
rect 9911 18244 9956 18272
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11977 18275 12035 18281
rect 11195 18244 11928 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11900 18216 11928 18244
rect 11977 18241 11989 18275
rect 12023 18272 12035 18275
rect 12621 18275 12679 18281
rect 12621 18272 12633 18275
rect 12023 18244 12633 18272
rect 12023 18241 12035 18244
rect 11977 18235 12035 18241
rect 12621 18241 12633 18244
rect 12667 18241 12679 18275
rect 12621 18235 12679 18241
rect 13538 18232 13544 18284
rect 13596 18272 13602 18284
rect 13633 18275 13691 18281
rect 13633 18272 13645 18275
rect 13596 18244 13645 18272
rect 13596 18232 13602 18244
rect 13633 18241 13645 18244
rect 13679 18272 13691 18275
rect 13722 18272 13728 18284
rect 13679 18244 13728 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 13722 18232 13728 18244
rect 13780 18272 13786 18284
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 13780 18244 14197 18272
rect 13780 18232 13786 18244
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 15286 18272 15292 18284
rect 15247 18244 15292 18272
rect 14185 18235 14243 18241
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 18380 18244 20269 18272
rect 18380 18232 18386 18244
rect 20257 18241 20269 18244
rect 20303 18272 20315 18275
rect 20346 18272 20352 18284
rect 20303 18244 20352 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 20824 18281 20852 18312
rect 20809 18275 20867 18281
rect 20809 18241 20821 18275
rect 20855 18272 20867 18275
rect 21266 18272 21272 18284
rect 20855 18244 21272 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 9548 18176 9593 18204
rect 9646 18176 11713 18204
rect 9548 18164 9554 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11882 18204 11888 18216
rect 11843 18176 11888 18204
rect 11701 18167 11759 18173
rect 3988 18108 4292 18136
rect 4338 18096 4344 18148
rect 4396 18136 4402 18148
rect 5261 18139 5319 18145
rect 5261 18136 5273 18139
rect 4396 18108 5273 18136
rect 4396 18096 4402 18108
rect 5261 18105 5273 18108
rect 5307 18105 5319 18139
rect 5261 18099 5319 18105
rect 5810 18096 5816 18148
rect 5868 18136 5874 18148
rect 8294 18136 8300 18148
rect 5868 18108 8300 18136
rect 5868 18096 5874 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 11716 18136 11744 18167
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18204 13231 18207
rect 14458 18204 14464 18216
rect 13219 18176 14464 18204
rect 13219 18173 13231 18176
rect 13173 18167 13231 18173
rect 13188 18136 13216 18167
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 17402 18204 17408 18216
rect 15611 18176 17408 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18204 18015 18207
rect 18003 18176 18920 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 11716 18108 13216 18136
rect 16761 18139 16819 18145
rect 16761 18105 16773 18139
rect 16807 18136 16819 18139
rect 16942 18136 16948 18148
rect 16807 18108 16948 18136
rect 16807 18105 16819 18108
rect 16761 18099 16819 18105
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 4430 18068 4436 18080
rect 2976 18040 4436 18068
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 4614 18068 4620 18080
rect 4575 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 6638 18068 6644 18080
rect 6599 18040 6644 18068
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 7374 18068 7380 18080
rect 7331 18040 7380 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 8478 18028 8484 18080
rect 8536 18068 8542 18080
rect 8941 18071 8999 18077
rect 8941 18068 8953 18071
rect 8536 18040 8953 18068
rect 8536 18028 8542 18040
rect 8941 18037 8953 18040
rect 8987 18037 8999 18071
rect 8941 18031 8999 18037
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10376 18040 10609 18068
rect 10376 18028 10382 18040
rect 10597 18037 10609 18040
rect 10643 18068 10655 18071
rect 10778 18068 10784 18080
rect 10643 18040 10784 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14792 18040 14933 18068
rect 14792 18028 14798 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 16206 18068 16212 18080
rect 16167 18040 16212 18068
rect 14921 18031 14979 18037
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 17221 18071 17279 18077
rect 17221 18068 17233 18071
rect 16356 18040 17233 18068
rect 16356 18028 16362 18040
rect 17221 18037 17233 18040
rect 17267 18068 17279 18071
rect 18230 18068 18236 18080
rect 17267 18040 18236 18068
rect 17267 18037 17279 18040
rect 17221 18031 17279 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 18506 18068 18512 18080
rect 18467 18040 18512 18068
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 18782 18068 18788 18080
rect 18743 18040 18788 18068
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18892 18068 18920 18176
rect 19058 18164 19064 18216
rect 19116 18204 19122 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 19116 18176 19257 18204
rect 19116 18164 19122 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 18966 18096 18972 18148
rect 19024 18136 19030 18148
rect 19352 18136 19380 18167
rect 19024 18108 19380 18136
rect 19024 18096 19030 18108
rect 19426 18068 19432 18080
rect 18892 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18068 19490 18080
rect 19797 18071 19855 18077
rect 19797 18068 19809 18071
rect 19484 18040 19809 18068
rect 19484 18028 19490 18040
rect 19797 18037 19809 18040
rect 19843 18037 19855 18071
rect 20438 18068 20444 18080
rect 20399 18040 20444 18068
rect 19797 18031 19855 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 1949 17867 2007 17873
rect 1949 17864 1961 17867
rect 1912 17836 1961 17864
rect 1912 17824 1918 17836
rect 1949 17833 1961 17836
rect 1995 17833 2007 17867
rect 1949 17827 2007 17833
rect 2593 17867 2651 17873
rect 2593 17833 2605 17867
rect 2639 17864 2651 17867
rect 2774 17864 2780 17876
rect 2639 17836 2780 17864
rect 2639 17833 2651 17836
rect 2593 17827 2651 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 5166 17824 5172 17876
rect 5224 17864 5230 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5224 17836 5641 17864
rect 5224 17824 5230 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 8754 17864 8760 17876
rect 6052 17836 8760 17864
rect 6052 17824 6058 17836
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 9585 17867 9643 17873
rect 9585 17864 9597 17867
rect 9456 17836 9597 17864
rect 9456 17824 9462 17836
rect 9585 17833 9597 17836
rect 9631 17833 9643 17867
rect 9585 17827 9643 17833
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 15194 17864 15200 17876
rect 9824 17836 15200 17864
rect 9824 17824 9830 17836
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 16117 17867 16175 17873
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 16482 17864 16488 17876
rect 16163 17836 16488 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 16577 17867 16635 17873
rect 16577 17833 16589 17867
rect 16623 17864 16635 17867
rect 17770 17864 17776 17876
rect 16623 17836 17776 17864
rect 16623 17833 16635 17836
rect 16577 17827 16635 17833
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 19116 17836 19257 17864
rect 19116 17824 19122 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 21266 17864 21272 17876
rect 19392 17836 20024 17864
rect 21227 17836 21272 17864
rect 19392 17824 19398 17836
rect 11054 17796 11060 17808
rect 6196 17768 11060 17796
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3292 17700 3801 17728
rect 3292 17688 3298 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 4798 17728 4804 17740
rect 4711 17700 4804 17728
rect 3789 17691 3847 17697
rect 4798 17688 4804 17700
rect 4856 17728 4862 17740
rect 6196 17728 6224 17768
rect 11054 17756 11060 17768
rect 11112 17756 11118 17808
rect 11517 17799 11575 17805
rect 11517 17765 11529 17799
rect 11563 17796 11575 17799
rect 12342 17796 12348 17808
rect 11563 17768 12348 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 12342 17756 12348 17768
rect 12400 17756 12406 17808
rect 16390 17756 16396 17808
rect 16448 17796 16454 17808
rect 17589 17799 17647 17805
rect 17589 17796 17601 17799
rect 16448 17768 17601 17796
rect 16448 17756 16454 17768
rect 17589 17765 17601 17768
rect 17635 17765 17647 17799
rect 17589 17759 17647 17765
rect 18064 17768 19840 17796
rect 4856 17700 6224 17728
rect 6273 17731 6331 17737
rect 4856 17688 4862 17700
rect 6273 17697 6285 17731
rect 6319 17697 6331 17731
rect 6914 17728 6920 17740
rect 6875 17700 6920 17728
rect 6273 17691 6331 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2406 17660 2412 17672
rect 2179 17632 2412 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17660 2835 17663
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 2823 17632 4261 17660
rect 2823 17629 2835 17632
rect 2777 17623 2835 17629
rect 4249 17629 4261 17632
rect 4295 17660 4307 17663
rect 6288 17660 6316 17691
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 9490 17728 9496 17740
rect 7975 17700 9496 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 10226 17728 10232 17740
rect 10187 17700 10232 17728
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 10686 17688 10692 17740
rect 10744 17728 10750 17740
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 10744 17700 12081 17728
rect 10744 17688 10750 17700
rect 12069 17697 12081 17700
rect 12115 17728 12127 17731
rect 12989 17731 13047 17737
rect 12989 17728 13001 17731
rect 12115 17700 13001 17728
rect 12115 17697 12127 17700
rect 12069 17691 12127 17697
rect 12989 17697 13001 17700
rect 13035 17697 13047 17731
rect 12989 17691 13047 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 18064 17728 18092 17768
rect 18230 17728 18236 17740
rect 15611 17700 18092 17728
rect 18191 17700 18236 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 19812 17737 19840 17768
rect 19797 17731 19855 17737
rect 18472 17700 19656 17728
rect 18472 17688 18478 17700
rect 6546 17660 6552 17672
rect 4295 17632 4844 17660
rect 6288 17632 6552 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4816 17604 4844 17632
rect 6546 17620 6552 17632
rect 6604 17660 6610 17672
rect 15838 17660 15844 17672
rect 6604 17632 15844 17660
rect 6604 17620 6610 17632
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16390 17660 16396 17672
rect 16351 17632 16396 17660
rect 16390 17620 16396 17632
rect 16448 17660 16454 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16448 17632 16957 17660
rect 16448 17620 16454 17632
rect 16945 17629 16957 17632
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18046 17660 18052 17672
rect 18003 17632 18052 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18046 17620 18052 17632
rect 18104 17620 18110 17672
rect 19628 17669 19656 17700
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 19886 17728 19892 17740
rect 19843 17700 19892 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 19996 17728 20024 17836
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 20809 17731 20867 17737
rect 20809 17728 20821 17731
rect 19996 17700 20821 17728
rect 20809 17697 20821 17700
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17629 19671 17663
rect 20714 17660 20720 17672
rect 19613 17623 19671 17629
rect 20640 17632 20720 17660
rect 4798 17552 4804 17604
rect 4856 17552 4862 17604
rect 4893 17595 4951 17601
rect 4893 17561 4905 17595
rect 4939 17592 4951 17595
rect 5718 17592 5724 17604
rect 4939 17564 5724 17592
rect 4939 17561 4951 17564
rect 4893 17555 4951 17561
rect 5718 17552 5724 17564
rect 5776 17552 5782 17604
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 8021 17595 8079 17601
rect 8021 17592 8033 17595
rect 7432 17564 8033 17592
rect 7432 17552 7438 17564
rect 8021 17561 8033 17564
rect 8067 17561 8079 17595
rect 8021 17555 8079 17561
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 8159 17564 8953 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8941 17561 8953 17564
rect 8987 17561 8999 17595
rect 8941 17555 8999 17561
rect 9398 17552 9404 17604
rect 9456 17592 9462 17604
rect 9766 17592 9772 17604
rect 9456 17564 9772 17592
rect 9456 17552 9462 17564
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 10045 17595 10103 17601
rect 10045 17561 10057 17595
rect 10091 17592 10103 17595
rect 10318 17592 10324 17604
rect 10091 17564 10324 17592
rect 10091 17561 10103 17564
rect 10045 17555 10103 17561
rect 10318 17552 10324 17564
rect 10376 17552 10382 17604
rect 10594 17552 10600 17604
rect 10652 17592 10658 17604
rect 11149 17595 11207 17601
rect 11149 17592 11161 17595
rect 10652 17564 11161 17592
rect 10652 17552 10658 17564
rect 11149 17561 11161 17564
rect 11195 17561 11207 17595
rect 11149 17555 11207 17561
rect 11885 17595 11943 17601
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 12529 17595 12587 17601
rect 12529 17592 12541 17595
rect 11931 17564 12541 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 12529 17561 12541 17564
rect 12575 17561 12587 17595
rect 12529 17555 12587 17561
rect 14274 17552 14280 17604
rect 14332 17592 14338 17604
rect 20640 17592 20668 17632
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 14332 17564 16528 17592
rect 14332 17552 14338 17564
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 1670 17524 1676 17536
rect 1627 17496 1676 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 3053 17527 3111 17533
rect 3053 17524 3065 17527
rect 3016 17496 3065 17524
rect 3016 17484 3022 17496
rect 3053 17493 3065 17496
rect 3099 17493 3111 17527
rect 3053 17487 3111 17493
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5040 17496 5085 17524
rect 5040 17484 5046 17496
rect 5166 17484 5172 17536
rect 5224 17524 5230 17536
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 5224 17496 5365 17524
rect 5224 17484 5230 17496
rect 5353 17493 5365 17496
rect 5399 17493 5411 17527
rect 5994 17524 6000 17536
rect 5955 17496 6000 17524
rect 5353 17487 5411 17493
rect 5994 17484 6000 17496
rect 6052 17484 6058 17536
rect 6089 17527 6147 17533
rect 6089 17493 6101 17527
rect 6135 17524 6147 17527
rect 6546 17524 6552 17536
rect 6135 17496 6552 17524
rect 6135 17493 6147 17496
rect 6089 17487 6147 17493
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7006 17524 7012 17536
rect 6696 17496 7012 17524
rect 6696 17484 6702 17496
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7466 17524 7472 17536
rect 7156 17496 7201 17524
rect 7427 17496 7472 17524
rect 7156 17484 7162 17496
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8444 17496 8493 17524
rect 8444 17484 8450 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 8481 17487 8539 17493
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9582 17524 9588 17536
rect 8812 17496 9588 17524
rect 8812 17484 8818 17496
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9732 17496 9965 17524
rect 9732 17484 9738 17496
rect 9953 17493 9965 17496
rect 9999 17493 10011 17527
rect 9953 17487 10011 17493
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10468 17496 10793 17524
rect 10468 17484 10474 17496
rect 10781 17493 10793 17496
rect 10827 17524 10839 17527
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 10827 17496 11989 17524
rect 10827 17493 10839 17496
rect 10781 17487 10839 17493
rect 11977 17493 11989 17496
rect 12023 17493 12035 17527
rect 11977 17487 12035 17493
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 13596 17496 15025 17524
rect 13596 17484 13602 17496
rect 15013 17493 15025 17496
rect 15059 17524 15071 17527
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15059 17496 15669 17524
rect 15059 17493 15071 17496
rect 15013 17487 15071 17493
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16500 17524 16528 17564
rect 19628 17564 20668 17592
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 15804 17496 15849 17524
rect 16500 17496 18061 17524
rect 15804 17484 15810 17496
rect 18049 17493 18061 17496
rect 18095 17524 18107 17527
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18095 17496 18613 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18601 17493 18613 17496
rect 18647 17524 18659 17527
rect 19628 17524 19656 17564
rect 18647 17496 19656 17524
rect 19705 17527 19763 17533
rect 18647 17493 18659 17496
rect 18601 17487 18659 17493
rect 19705 17493 19717 17527
rect 19751 17524 19763 17527
rect 19978 17524 19984 17536
rect 19751 17496 19984 17524
rect 19751 17493 19763 17496
rect 19705 17487 19763 17493
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 20438 17524 20444 17536
rect 20303 17496 20444 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20622 17524 20628 17536
rect 20583 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 20898 17524 20904 17536
rect 20763 17496 20904 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1486 17320 1492 17332
rect 1447 17292 1492 17320
rect 1486 17280 1492 17292
rect 1544 17280 1550 17332
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 4062 17320 4068 17332
rect 3936 17292 4068 17320
rect 3936 17280 3942 17292
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4212 17292 4445 17320
rect 4212 17280 4218 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 5166 17320 5172 17332
rect 5127 17292 5172 17320
rect 4433 17283 4491 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 5810 17280 5816 17332
rect 5868 17320 5874 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 5868 17292 6837 17320
rect 5868 17280 5874 17292
rect 6825 17289 6837 17292
rect 6871 17320 6883 17323
rect 8386 17320 8392 17332
rect 6871 17292 8064 17320
rect 8347 17292 8392 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 3326 17212 3332 17264
rect 3384 17252 3390 17264
rect 3973 17255 4031 17261
rect 3973 17252 3985 17255
rect 3384 17224 3985 17252
rect 3384 17212 3390 17224
rect 3973 17221 3985 17224
rect 4019 17221 4031 17255
rect 3973 17215 4031 17221
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 5077 17255 5135 17261
rect 5077 17252 5089 17255
rect 4672 17224 5089 17252
rect 4672 17212 4678 17224
rect 5077 17221 5089 17224
rect 5123 17221 5135 17255
rect 5077 17215 5135 17221
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 2958 17184 2964 17196
rect 2919 17156 2964 17184
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17184 3479 17187
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3467 17156 4077 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 6917 17187 6975 17193
rect 4065 17147 4123 17153
rect 4540 17156 6868 17184
rect 1578 17008 1584 17060
rect 1636 17048 1642 17060
rect 3436 17048 3464 17147
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17116 3939 17119
rect 4430 17116 4436 17128
rect 3927 17088 4436 17116
rect 3927 17085 3939 17088
rect 3881 17079 3939 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 1636 17020 3464 17048
rect 1636 17008 1642 17020
rect 2130 16980 2136 16992
rect 2091 16952 2136 16980
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 2866 16980 2872 16992
rect 2823 16952 2872 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 4540 16980 4568 17156
rect 5350 17116 5356 17128
rect 5311 17088 5356 17116
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17085 6791 17119
rect 6840 17116 6868 17156
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 6963 17156 7573 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 8036 17184 8064 17292
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 8536 17292 8581 17320
rect 8536 17280 8542 17292
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8720 17292 9045 17320
rect 8720 17280 8726 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9950 17320 9956 17332
rect 9033 17283 9091 17289
rect 9232 17292 9956 17320
rect 9232 17184 9260 17292
rect 9950 17280 9956 17292
rect 10008 17320 10014 17332
rect 10410 17320 10416 17332
rect 10008 17292 10416 17320
rect 10008 17280 10014 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 10594 17280 10600 17332
rect 10652 17320 10658 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10652 17292 10701 17320
rect 10652 17280 10658 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 14274 17320 14280 17332
rect 10689 17283 10747 17289
rect 12406 17292 13768 17320
rect 14235 17292 14280 17320
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 12406 17252 12434 17292
rect 9640 17224 12434 17252
rect 9640 17212 9646 17224
rect 9398 17184 9404 17196
rect 8036 17156 9260 17184
rect 9359 17156 9404 17184
rect 7561 17147 7619 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10060 17156 10793 17184
rect 8662 17116 8668 17128
rect 6840 17088 8340 17116
rect 8623 17088 8668 17116
rect 6733 17079 6791 17085
rect 6748 17048 6776 17079
rect 7834 17048 7840 17060
rect 6748 17020 7840 17048
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 4706 16980 4712 16992
rect 3108 16952 4568 16980
rect 4667 16952 4712 16980
rect 3108 16940 3114 16952
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 5810 16940 5816 16992
rect 5868 16980 5874 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5868 16952 5917 16980
rect 5868 16940 5874 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 7282 16980 7288 16992
rect 7243 16952 7288 16980
rect 5905 16943 5963 16949
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 8018 16980 8024 16992
rect 7979 16952 8024 16980
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 8312 16980 8340 17088
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 9508 17048 9536 17079
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 9640 17088 9685 17116
rect 9640 17076 9646 17088
rect 8444 17020 9536 17048
rect 8444 17008 8450 17020
rect 10060 16989 10088 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12023 17156 12633 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 13740 17184 13768 17292
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15286 17320 15292 17332
rect 14783 17292 15292 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15838 17280 15844 17332
rect 15896 17320 15902 17332
rect 16850 17320 16856 17332
rect 15896 17292 16856 17320
rect 15896 17280 15902 17292
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 18690 17280 18696 17332
rect 18748 17320 18754 17332
rect 20806 17320 20812 17332
rect 18748 17292 19932 17320
rect 20767 17292 20812 17320
rect 18748 17280 18754 17292
rect 13814 17212 13820 17264
rect 13872 17252 13878 17264
rect 18046 17252 18052 17264
rect 13872 17224 18052 17252
rect 13872 17212 13878 17224
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 19794 17252 19800 17264
rect 19755 17224 19800 17252
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 19904 17252 19932 17292
rect 20806 17280 20812 17292
rect 20864 17280 20870 17332
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 19904 17224 20729 17252
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20717 17215 20775 17221
rect 14369 17187 14427 17193
rect 13740 17156 14320 17184
rect 12621 17147 12679 17153
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 10597 17079 10655 17085
rect 10612 17048 10640 17079
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 14185 17119 14243 17125
rect 11940 17088 11985 17116
rect 11940 17076 11946 17088
rect 14185 17085 14197 17119
rect 14231 17085 14243 17119
rect 14292 17116 14320 17156
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 15013 17187 15071 17193
rect 15013 17184 15025 17187
rect 14415 17156 15025 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 15013 17153 15025 17156
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16942 17184 16948 17196
rect 16715 17156 16948 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16942 17144 16948 17156
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 20070 17184 20076 17196
rect 20031 17156 20076 17184
rect 17221 17147 17279 17153
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 18046 17116 18052 17128
rect 14292 17088 18052 17116
rect 14185 17079 14243 17085
rect 11808 17048 11836 17076
rect 10612 17020 11836 17048
rect 14200 17048 14228 17079
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 20806 17076 20812 17128
rect 20864 17116 20870 17128
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20864 17088 20913 17116
rect 20864 17076 20870 17088
rect 20901 17085 20913 17088
rect 20947 17085 20959 17119
rect 20901 17079 20959 17085
rect 15378 17048 15384 17060
rect 14200 17020 15384 17048
rect 15378 17008 15384 17020
rect 15436 17048 15442 17060
rect 16114 17048 16120 17060
rect 15436 17020 16120 17048
rect 15436 17008 15442 17020
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 16853 17051 16911 17057
rect 16853 17017 16865 17051
rect 16899 17048 16911 17051
rect 17954 17048 17960 17060
rect 16899 17020 17960 17048
rect 16899 17017 16911 17020
rect 16853 17011 16911 17017
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 10045 16983 10103 16989
rect 10045 16980 10057 16983
rect 8312 16952 10057 16980
rect 10045 16949 10057 16952
rect 10091 16949 10103 16983
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 10045 16943 10103 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 12986 16980 12992 16992
rect 12391 16952 12992 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 13320 16952 13645 16980
rect 13320 16940 13326 16952
rect 13633 16949 13645 16952
rect 13679 16980 13691 16983
rect 14274 16980 14280 16992
rect 13679 16952 14280 16980
rect 13679 16949 13691 16952
rect 13633 16943 13691 16949
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 17589 16983 17647 16989
rect 17589 16980 17601 16983
rect 17000 16952 17601 16980
rect 17000 16940 17006 16952
rect 17589 16949 17601 16952
rect 17635 16949 17647 16983
rect 17589 16943 17647 16949
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 18598 16980 18604 16992
rect 18555 16952 18604 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 3326 16776 3332 16788
rect 1728 16748 2774 16776
rect 3287 16748 3332 16776
rect 1728 16736 1734 16748
rect 2746 16708 2774 16748
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 5810 16776 5816 16788
rect 3936 16748 5816 16776
rect 3936 16736 3942 16748
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7190 16776 7196 16788
rect 6972 16748 7196 16776
rect 6972 16736 6978 16748
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8444 16748 9137 16776
rect 8444 16736 8450 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 15654 16776 15660 16788
rect 9125 16739 9183 16745
rect 11072 16748 15660 16776
rect 4522 16708 4528 16720
rect 2746 16680 4292 16708
rect 4483 16680 4528 16708
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16640 4031 16643
rect 4154 16640 4160 16652
rect 4019 16612 4160 16640
rect 4019 16609 4031 16612
rect 3973 16603 4031 16609
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4264 16640 4292 16680
rect 4522 16668 4528 16680
rect 4580 16668 4586 16720
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 6181 16711 6239 16717
rect 6181 16708 6193 16711
rect 5500 16680 6193 16708
rect 5500 16668 5506 16680
rect 6181 16677 6193 16680
rect 6227 16708 6239 16711
rect 7098 16708 7104 16720
rect 6227 16680 7104 16708
rect 6227 16677 6239 16680
rect 6181 16671 6239 16677
rect 7098 16668 7104 16680
rect 7156 16708 7162 16720
rect 8294 16708 8300 16720
rect 7156 16680 8300 16708
rect 7156 16668 7162 16680
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8573 16711 8631 16717
rect 8573 16677 8585 16711
rect 8619 16708 8631 16711
rect 8754 16708 8760 16720
rect 8619 16680 8760 16708
rect 8619 16677 8631 16680
rect 8573 16671 8631 16677
rect 8754 16668 8760 16680
rect 8812 16708 8818 16720
rect 9398 16708 9404 16720
rect 8812 16680 9404 16708
rect 8812 16668 8818 16680
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 6549 16643 6607 16649
rect 4264 16612 6500 16640
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2961 16575 3019 16581
rect 2271 16544 2912 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2038 16464 2044 16516
rect 2096 16504 2102 16516
rect 2685 16507 2743 16513
rect 2685 16504 2697 16507
rect 2096 16476 2697 16504
rect 2096 16464 2102 16476
rect 2685 16473 2697 16476
rect 2731 16473 2743 16507
rect 2884 16504 2912 16544
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 4706 16572 4712 16584
rect 3007 16544 4712 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 6472 16572 6500 16612
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 7006 16640 7012 16652
rect 6595 16612 7012 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 7006 16600 7012 16612
rect 7064 16640 7070 16652
rect 7374 16640 7380 16652
rect 7064 16612 7380 16640
rect 7064 16600 7070 16612
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 7926 16600 7932 16652
rect 7984 16640 7990 16652
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 7984 16612 9505 16640
rect 7984 16600 7990 16612
rect 9493 16609 9505 16612
rect 9539 16640 9551 16643
rect 10045 16643 10103 16649
rect 9539 16612 9720 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 6472 16544 6776 16572
rect 3418 16504 3424 16516
rect 2884 16476 3424 16504
rect 2685 16467 2743 16473
rect 3418 16464 3424 16476
rect 3476 16464 3482 16516
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16504 4123 16507
rect 4338 16504 4344 16516
rect 4111 16476 4344 16504
rect 4111 16473 4123 16476
rect 4065 16467 4123 16473
rect 4338 16464 4344 16476
rect 4396 16464 4402 16516
rect 5350 16504 5356 16516
rect 4448 16476 5356 16504
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 4448 16436 4476 16476
rect 5350 16464 5356 16476
rect 5408 16464 5414 16516
rect 5810 16504 5816 16516
rect 5723 16476 5816 16504
rect 5810 16464 5816 16476
rect 5868 16504 5874 16516
rect 6638 16504 6644 16516
rect 5868 16476 6644 16504
rect 5868 16464 5874 16476
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 6748 16504 6776 16544
rect 6914 16532 6920 16584
rect 6972 16572 6978 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 6972 16544 8125 16572
rect 6972 16532 6978 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 9692 16572 9720 16612
rect 10045 16609 10057 16643
rect 10091 16640 10103 16643
rect 10962 16640 10968 16652
rect 10091 16612 10968 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11072 16649 11100 16748
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 16209 16779 16267 16785
rect 16209 16776 16221 16779
rect 15804 16748 16221 16776
rect 15804 16736 15810 16748
rect 16209 16745 16221 16748
rect 16255 16745 16267 16779
rect 16209 16739 16267 16745
rect 19981 16779 20039 16785
rect 19981 16745 19993 16779
rect 20027 16776 20039 16779
rect 20070 16776 20076 16788
rect 20027 16748 20076 16776
rect 20027 16745 20039 16748
rect 19981 16739 20039 16745
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 11146 16668 11152 16720
rect 11204 16708 11210 16720
rect 21082 16708 21088 16720
rect 11204 16680 12940 16708
rect 11204 16668 11210 16680
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11882 16640 11888 16652
rect 11843 16612 11888 16640
rect 11057 16603 11115 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 12912 16649 12940 16680
rect 16960 16680 21088 16708
rect 16960 16652 16988 16680
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15841 16643 15899 16649
rect 15841 16640 15853 16643
rect 15528 16612 15853 16640
rect 15528 16600 15534 16612
rect 15841 16609 15853 16612
rect 15887 16640 15899 16643
rect 16390 16640 16396 16652
rect 15887 16612 16396 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16390 16600 16396 16612
rect 16448 16640 16454 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16448 16612 16681 16640
rect 16448 16600 16454 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 16669 16603 16727 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 16942 16640 16948 16652
rect 16899 16612 16948 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 17092 16612 17785 16640
rect 17092 16600 17098 16612
rect 17773 16609 17785 16612
rect 17819 16609 17831 16643
rect 20438 16640 20444 16652
rect 20399 16612 20444 16640
rect 17773 16603 17831 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 20588 16612 20633 16640
rect 20588 16600 20594 16612
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 9692 16544 10241 16572
rect 8113 16535 8171 16541
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 11238 16572 11244 16584
rect 11199 16544 11244 16572
rect 10229 16535 10287 16541
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12986 16572 12992 16584
rect 12947 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 18598 16572 18604 16584
rect 17635 16544 18604 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 18782 16572 18788 16584
rect 18743 16544 18788 16572
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20680 16544 21005 16572
rect 20680 16532 20686 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 6748 16476 6960 16504
rect 4890 16436 4896 16448
rect 4203 16408 4476 16436
rect 4851 16408 4896 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 5132 16408 5273 16436
rect 5132 16396 5138 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 5718 16396 5724 16448
rect 5776 16436 5782 16448
rect 6822 16436 6828 16448
rect 5776 16408 6828 16436
rect 5776 16396 5782 16408
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6932 16445 6960 16476
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 7745 16507 7803 16513
rect 7745 16504 7757 16507
rect 7156 16476 7757 16504
rect 7156 16464 7162 16476
rect 7745 16473 7757 16476
rect 7791 16473 7803 16507
rect 15562 16504 15568 16516
rect 7745 16467 7803 16473
rect 11624 16476 15568 16504
rect 6917 16439 6975 16445
rect 6917 16405 6929 16439
rect 6963 16436 6975 16439
rect 7006 16436 7012 16448
rect 6963 16408 7012 16436
rect 6963 16405 6975 16408
rect 6917 16399 6975 16405
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 10134 16436 10140 16448
rect 10095 16408 10140 16436
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 11624 16445 11652 16476
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 17681 16507 17739 16513
rect 16080 16476 17264 16504
rect 16080 16464 16086 16476
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 10643 16408 11161 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16405 11667 16439
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 11609 16399 11667 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 17236 16445 17264 16476
rect 17681 16473 17693 16507
rect 17727 16504 17739 16507
rect 17954 16504 17960 16516
rect 17727 16476 17960 16504
rect 17727 16473 17739 16476
rect 17681 16467 17739 16473
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 18509 16507 18567 16513
rect 18509 16473 18521 16507
rect 18555 16504 18567 16507
rect 20714 16504 20720 16516
rect 18555 16476 20720 16504
rect 18555 16473 18567 16476
rect 18509 16467 18567 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 16577 16439 16635 16445
rect 16577 16436 16589 16439
rect 16448 16408 16589 16436
rect 16448 16396 16454 16408
rect 16577 16405 16589 16408
rect 16623 16405 16635 16439
rect 16577 16399 16635 16405
rect 17221 16439 17279 16445
rect 17221 16405 17233 16439
rect 17267 16405 17279 16439
rect 17221 16399 17279 16405
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 18104 16408 20361 16436
rect 18104 16396 18110 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 21174 16436 21180 16448
rect 21135 16408 21180 16436
rect 20349 16399 20407 16405
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2774 16232 2780 16244
rect 2455 16204 2780 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5077 16235 5135 16241
rect 5077 16232 5089 16235
rect 5040 16204 5089 16232
rect 5040 16192 5046 16204
rect 5077 16201 5089 16204
rect 5123 16201 5135 16235
rect 5077 16195 5135 16201
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 5810 16232 5816 16244
rect 5491 16204 5816 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 6880 16204 7573 16232
rect 6880 16192 6886 16204
rect 7561 16201 7573 16204
rect 7607 16201 7619 16235
rect 7561 16195 7619 16201
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 9766 16232 9772 16244
rect 7708 16204 9772 16232
rect 7708 16192 7714 16204
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 7006 16164 7012 16176
rect 4028 16136 6776 16164
rect 6919 16136 7012 16164
rect 4028 16124 4034 16136
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 4430 16096 4436 16108
rect 2639 16068 3004 16096
rect 4391 16068 4436 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 2976 15969 3004 16068
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 4614 16056 4620 16108
rect 4672 16096 4678 16108
rect 4672 16068 5396 16096
rect 4672 16056 4678 16068
rect 4522 16028 4528 16040
rect 4483 16000 4528 16028
rect 4522 15988 4528 16000
rect 4580 15988 4586 16040
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 16028 4767 16031
rect 4890 16028 4896 16040
rect 4755 16000 4896 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 4890 15988 4896 16000
rect 4948 16028 4954 16040
rect 5258 16028 5264 16040
rect 4948 16000 5264 16028
rect 4948 15988 4954 16000
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 5368 16028 5396 16068
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5500 16068 5549 16096
rect 5500 16056 5506 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 5721 16031 5779 16037
rect 5721 16028 5733 16031
rect 5368 16000 5733 16028
rect 5721 15997 5733 16000
rect 5767 16028 5779 16031
rect 5767 16000 6684 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 2961 15963 3019 15969
rect 2961 15929 2973 15963
rect 3007 15960 3019 15963
rect 5810 15960 5816 15972
rect 3007 15932 5816 15960
rect 3007 15929 3019 15932
rect 2961 15923 3019 15929
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1857 15895 1915 15901
rect 1857 15892 1869 15895
rect 1452 15864 1869 15892
rect 1452 15852 1458 15864
rect 1857 15861 1869 15864
rect 1903 15861 1915 15895
rect 1857 15855 1915 15861
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 4338 15892 4344 15904
rect 4111 15864 4344 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 6656 15892 6684 16000
rect 6748 15960 6776 16136
rect 7006 16124 7012 16136
rect 7064 16164 7070 16176
rect 8110 16164 8116 16176
rect 7064 16136 8116 16164
rect 7064 16124 7070 16136
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 6914 16096 6920 16108
rect 6875 16068 6920 16096
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7432 16068 7941 16096
rect 7432 16056 7438 16068
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 8018 16028 8024 16040
rect 7156 16000 7201 16028
rect 7979 16000 8024 16028
rect 7156 15988 7162 16000
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8312 16028 8340 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10192 16204 11529 16232
rect 10192 16192 10198 16204
rect 11517 16201 11529 16204
rect 11563 16232 11575 16235
rect 12066 16232 12072 16244
rect 11563 16204 12072 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 13722 16232 13728 16244
rect 13504 16204 13728 16232
rect 13504 16192 13510 16204
rect 13722 16192 13728 16204
rect 13780 16232 13786 16244
rect 14185 16235 14243 16241
rect 14185 16232 14197 16235
rect 13780 16204 14197 16232
rect 13780 16192 13786 16204
rect 14185 16201 14197 16204
rect 14231 16201 14243 16235
rect 14185 16195 14243 16201
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16448 16204 16773 16232
rect 16448 16192 16454 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 17727 16204 18337 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18325 16195 18383 16201
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18564 16204 18797 16232
rect 18564 16192 18570 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 8662 16124 8668 16176
rect 8720 16164 8726 16176
rect 10238 16167 10296 16173
rect 10238 16164 10250 16167
rect 8720 16136 10250 16164
rect 8720 16124 8726 16136
rect 10238 16133 10250 16136
rect 10284 16164 10296 16167
rect 19058 16164 19064 16176
rect 10284 16136 12434 16164
rect 10284 16133 10296 16136
rect 10238 16127 10296 16133
rect 10594 16096 10600 16108
rect 8251 16000 8340 16028
rect 8680 16068 10600 16096
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 6748 15932 8064 15960
rect 7650 15892 7656 15904
rect 6656 15864 7656 15892
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 8036 15892 8064 15932
rect 8202 15892 8208 15904
rect 8036 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15892 8266 15904
rect 8680 15901 8708 16068
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 12406 16096 12434 16136
rect 17604 16136 19064 16164
rect 13722 16096 13728 16108
rect 12406 16068 13728 16096
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 17604 16096 17632 16136
rect 19058 16124 19064 16136
rect 19116 16124 19122 16176
rect 20622 16164 20628 16176
rect 20583 16136 20628 16164
rect 20622 16124 20628 16136
rect 20680 16124 20686 16176
rect 14016 16068 14964 16096
rect 14016 16037 14044 16068
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 14001 16031 14059 16037
rect 10551 16000 10824 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 10796 15904 10824 16000
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 14108 15960 14136 15991
rect 13464 15932 14136 15960
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8260 15864 8677 15892
rect 8260 15852 8266 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 9125 15895 9183 15901
rect 9125 15861 9137 15895
rect 9171 15892 9183 15895
rect 9398 15892 9404 15904
rect 9171 15864 9404 15892
rect 9171 15861 9183 15864
rect 9125 15855 9183 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 13464 15901 13492 15932
rect 14936 15901 14964 16068
rect 17512 16068 17632 16096
rect 17512 16037 17540 16068
rect 18506 16056 18512 16108
rect 18564 16096 18570 16108
rect 18693 16099 18751 16105
rect 18693 16096 18705 16099
rect 18564 16068 18705 16096
rect 18564 16056 18570 16068
rect 18693 16065 18705 16068
rect 18739 16065 18751 16099
rect 20346 16096 20352 16108
rect 20307 16068 20352 16096
rect 18693 16059 18751 16065
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 17589 16031 17647 16037
rect 17589 15997 17601 16031
rect 17635 16028 17647 16031
rect 17770 16028 17776 16040
rect 17635 16000 17776 16028
rect 17635 15997 17647 16000
rect 17589 15991 17647 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 16028 19027 16031
rect 19794 16028 19800 16040
rect 19015 16000 19800 16028
rect 19015 15997 19027 16000
rect 18969 15991 19027 15997
rect 19794 15988 19800 16000
rect 19852 15988 19858 16040
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19944 16000 19993 16028
rect 19944 15988 19950 16000
rect 19981 15997 19993 16000
rect 20027 16028 20039 16031
rect 21100 16028 21128 16059
rect 20027 16000 21128 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 18046 15960 18052 15972
rect 18007 15932 18052 15960
rect 18046 15920 18052 15932
rect 18104 15920 18110 15972
rect 21266 15960 21272 15972
rect 21227 15932 21272 15960
rect 21266 15920 21272 15932
rect 21324 15920 21330 15972
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13136 15864 13461 15892
rect 13136 15852 13142 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 16114 15892 16120 15904
rect 14967 15864 16120 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 16114 15852 16120 15864
rect 16172 15892 16178 15904
rect 16298 15892 16304 15904
rect 16172 15864 16304 15892
rect 16172 15852 16178 15864
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 19518 15852 19524 15904
rect 19576 15892 19582 15904
rect 19886 15892 19892 15904
rect 19576 15864 19892 15892
rect 19576 15852 19582 15864
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 4430 15688 4436 15700
rect 4391 15660 4436 15688
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 8018 15648 8024 15700
rect 8076 15688 8082 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 8076 15660 8217 15688
rect 8076 15648 8082 15660
rect 8205 15657 8217 15660
rect 8251 15657 8263 15691
rect 8205 15651 8263 15657
rect 9232 15660 10180 15688
rect 2314 15620 2320 15632
rect 2275 15592 2320 15620
rect 2314 15580 2320 15592
rect 2372 15580 2378 15632
rect 6917 15623 6975 15629
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 9232 15620 9260 15660
rect 6963 15592 9260 15620
rect 10152 15620 10180 15660
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 10284 15660 10609 15688
rect 10284 15648 10290 15660
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 10597 15651 10655 15657
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 13633 15691 13691 15697
rect 13633 15688 13645 15691
rect 13504 15660 13645 15688
rect 13504 15648 13510 15660
rect 13633 15657 13645 15660
rect 13679 15657 13691 15691
rect 16298 15688 16304 15700
rect 13633 15651 13691 15657
rect 14384 15660 16304 15688
rect 11698 15620 11704 15632
rect 10152 15592 11704 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 14384 15620 14412 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16942 15688 16948 15700
rect 16903 15660 16948 15688
rect 16942 15648 16948 15660
rect 17000 15688 17006 15700
rect 17218 15688 17224 15700
rect 17000 15660 17224 15688
rect 17000 15648 17006 15660
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 19981 15691 20039 15697
rect 19981 15688 19993 15691
rect 19306 15660 19993 15688
rect 19306 15620 19334 15660
rect 19981 15657 19993 15660
rect 20027 15688 20039 15691
rect 20346 15688 20352 15700
rect 20027 15660 20352 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 12406 15592 14412 15620
rect 16592 15592 19334 15620
rect 5074 15552 5080 15564
rect 5035 15524 5080 15552
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15552 6423 15555
rect 7190 15552 7196 15564
rect 6411 15524 7196 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 7650 15552 7656 15564
rect 7611 15524 7656 15552
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8754 15552 8760 15564
rect 8536 15524 8760 15552
rect 8536 15512 8542 15524
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 12406 15552 12434 15592
rect 16592 15552 16620 15592
rect 18506 15552 18512 15564
rect 10652 15524 12434 15552
rect 16500 15524 16620 15552
rect 18467 15524 18512 15552
rect 10652 15512 10658 15524
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 3329 15487 3387 15493
rect 3329 15484 3341 15487
rect 2547 15456 3341 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 3329 15453 3341 15456
rect 3375 15484 3387 15487
rect 4614 15484 4620 15496
rect 3375 15456 4620 15484
rect 3375 15453 3387 15456
rect 3329 15447 3387 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 6546 15484 6552 15496
rect 4724 15456 5580 15484
rect 6507 15456 6552 15484
rect 3050 15376 3056 15428
rect 3108 15416 3114 15428
rect 4724 15416 4752 15456
rect 3108 15388 4752 15416
rect 4801 15419 4859 15425
rect 3108 15376 3114 15388
rect 4801 15385 4813 15419
rect 4847 15416 4859 15419
rect 5445 15419 5503 15425
rect 5445 15416 5457 15419
rect 4847 15388 5457 15416
rect 4847 15385 4859 15388
rect 4801 15379 4859 15385
rect 5445 15385 5457 15388
rect 5491 15385 5503 15419
rect 5445 15379 5503 15385
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2924 15320 2973 15348
rect 2924 15308 2930 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 2961 15311 3019 15317
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 4157 15351 4215 15357
rect 4157 15348 4169 15351
rect 3292 15320 4169 15348
rect 3292 15308 3298 15320
rect 4157 15317 4169 15320
rect 4203 15348 4215 15351
rect 4893 15351 4951 15357
rect 4893 15348 4905 15351
rect 4203 15320 4905 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 4893 15317 4905 15320
rect 4939 15317 4951 15351
rect 5552 15348 5580 15456
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 9214 15484 9220 15496
rect 6748 15456 8616 15484
rect 9175 15456 9220 15484
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 6638 15416 6644 15428
rect 6503 15388 6644 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 6638 15376 6644 15388
rect 6696 15376 6702 15428
rect 6748 15348 6776 15456
rect 8481 15419 8539 15425
rect 8481 15416 8493 15419
rect 7760 15388 8493 15416
rect 7760 15360 7788 15388
rect 8481 15385 8493 15388
rect 8527 15385 8539 15419
rect 8481 15379 8539 15385
rect 7742 15348 7748 15360
rect 5552 15320 6776 15348
rect 7703 15320 7748 15348
rect 4893 15311 4951 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 8202 15348 8208 15360
rect 7883 15320 8208 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8588 15348 8616 15456
rect 9214 15444 9220 15456
rect 9272 15484 9278 15496
rect 10778 15484 10784 15496
rect 9272 15456 10784 15484
rect 9272 15444 9278 15456
rect 10778 15444 10784 15456
rect 10836 15484 10842 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 10836 15456 10885 15484
rect 10836 15444 10842 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 13262 15484 13268 15496
rect 10873 15447 10931 15453
rect 12406 15456 13268 15484
rect 9306 15376 9312 15428
rect 9364 15416 9370 15428
rect 9462 15419 9520 15425
rect 9462 15416 9474 15419
rect 9364 15388 9474 15416
rect 9364 15376 9370 15388
rect 9462 15385 9474 15388
rect 9508 15416 9520 15419
rect 10962 15416 10968 15428
rect 9508 15388 10968 15416
rect 9508 15385 9520 15388
rect 9462 15379 9520 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 12406 15348 12434 15456
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 16500 15484 16528 15524
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 14516 15456 16528 15484
rect 16577 15487 16635 15493
rect 14516 15444 14522 15456
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16942 15484 16948 15496
rect 16623 15456 16948 15484
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16942 15444 16948 15456
rect 17000 15484 17006 15496
rect 20714 15484 20720 15496
rect 17000 15456 17356 15484
rect 20675 15456 20720 15484
rect 17000 15444 17006 15456
rect 16332 15419 16390 15425
rect 16332 15385 16344 15419
rect 16378 15416 16390 15419
rect 17034 15416 17040 15428
rect 16378 15388 17040 15416
rect 16378 15385 16390 15388
rect 16332 15379 16390 15385
rect 17034 15376 17040 15388
rect 17092 15376 17098 15428
rect 8588 15320 12434 15348
rect 15197 15351 15255 15357
rect 15197 15317 15209 15351
rect 15243 15348 15255 15351
rect 15378 15348 15384 15360
rect 15243 15320 15384 15348
rect 15243 15317 15255 15320
rect 15197 15311 15255 15317
rect 15378 15308 15384 15320
rect 15436 15348 15442 15360
rect 15838 15348 15844 15360
rect 15436 15320 15844 15348
rect 15436 15308 15442 15320
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 17328 15357 17356 15456
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 20349 15419 20407 15425
rect 20349 15385 20361 15419
rect 20395 15385 20407 15419
rect 20349 15379 20407 15385
rect 17313 15351 17371 15357
rect 17313 15317 17325 15351
rect 17359 15348 17371 15351
rect 18322 15348 18328 15360
rect 17359 15320 18328 15348
rect 17359 15317 17371 15320
rect 17313 15311 17371 15317
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19576 15320 19625 15348
rect 19576 15308 19582 15320
rect 19613 15317 19625 15320
rect 19659 15348 19671 15351
rect 20364 15348 20392 15379
rect 19659 15320 20392 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 20901 15351 20959 15357
rect 20901 15348 20913 15351
rect 20496 15320 20913 15348
rect 20496 15308 20502 15320
rect 20901 15317 20913 15320
rect 20947 15317 20959 15351
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 20901 15311 20959 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 3326 15104 3332 15156
rect 3384 15144 3390 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3384 15116 3893 15144
rect 3384 15104 3390 15116
rect 3881 15113 3893 15116
rect 3927 15144 3939 15147
rect 4062 15144 4068 15156
rect 3927 15116 4068 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 5500 15116 8616 15144
rect 5500 15104 5506 15116
rect 2406 15036 2412 15088
rect 2464 15076 2470 15088
rect 7745 15079 7803 15085
rect 7745 15076 7757 15079
rect 2464 15048 7757 15076
rect 2464 15036 2470 15048
rect 7745 15045 7757 15048
rect 7791 15076 7803 15079
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 7791 15048 8309 15076
rect 7791 15045 7803 15048
rect 7745 15039 7803 15045
rect 8297 15045 8309 15048
rect 8343 15076 8355 15079
rect 8478 15076 8484 15088
rect 8343 15048 8484 15076
rect 8343 15045 8355 15048
rect 8297 15039 8355 15045
rect 8478 15036 8484 15048
rect 8536 15036 8542 15088
rect 8588 15076 8616 15116
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 13262 15144 13268 15156
rect 8812 15116 13268 15144
rect 8812 15104 8818 15116
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 14826 15144 14832 15156
rect 13372 15116 14688 15144
rect 14787 15116 14832 15144
rect 13372 15076 13400 15116
rect 8588 15048 13400 15076
rect 14660 15076 14688 15116
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15930 15144 15936 15156
rect 15580 15116 15936 15144
rect 15470 15076 15476 15088
rect 14660 15048 15476 15076
rect 15470 15036 15476 15048
rect 15528 15036 15534 15088
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 2866 15008 2872 15020
rect 2827 14980 2872 15008
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 14977 3203 15011
rect 4982 15008 4988 15020
rect 4943 14980 4988 15008
rect 3145 14971 3203 14977
rect 2133 14943 2191 14949
rect 2133 14909 2145 14943
rect 2179 14940 2191 14943
rect 3160 14940 3188 14971
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5994 15008 6000 15020
rect 5123 14980 6000 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 5258 14940 5264 14952
rect 2179 14912 3188 14940
rect 5219 14912 5264 14940
rect 2179 14909 2191 14912
rect 2133 14903 2191 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5592 14912 5917 14940
rect 5592 14900 5598 14912
rect 5905 14909 5917 14912
rect 5951 14940 5963 14943
rect 6546 14940 6552 14952
rect 5951 14912 6552 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 4706 14832 4712 14884
rect 4764 14872 4770 14884
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 4764 14844 6929 14872
rect 4764 14832 4770 14844
rect 6917 14841 6929 14844
rect 6963 14872 6975 14875
rect 7668 14872 7696 14971
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9272 14980 9689 15008
rect 9272 14968 9278 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9944 15011 10002 15017
rect 9944 15008 9956 15011
rect 9824 14980 9956 15008
rect 9824 14968 9830 14980
rect 9944 14977 9956 14980
rect 9990 15008 10002 15011
rect 10410 15008 10416 15020
rect 9990 14980 10416 15008
rect 9990 14977 10002 14980
rect 9944 14971 10002 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13538 15008 13544 15020
rect 13495 14980 13544 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 13716 15011 13774 15017
rect 13716 14977 13728 15011
rect 13762 15008 13774 15011
rect 15580 15008 15608 15116
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 16942 15104 16948 15156
rect 17000 15104 17006 15156
rect 16960 15076 16988 15104
rect 16684 15048 16988 15076
rect 16684 15017 16712 15048
rect 18690 15036 18696 15088
rect 18748 15076 18754 15088
rect 20134 15079 20192 15085
rect 20134 15076 20146 15079
rect 18748 15048 20146 15076
rect 18748 15036 18754 15048
rect 20134 15045 20146 15048
rect 20180 15045 20192 15079
rect 20134 15039 20192 15045
rect 13762 14980 15608 15008
rect 16669 15011 16727 15017
rect 13762 14977 13774 14980
rect 13716 14971 13774 14977
rect 16669 14977 16681 15011
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16936 15011 16994 15017
rect 16936 14977 16948 15011
rect 16982 15008 16994 15011
rect 17218 15008 17224 15020
rect 16982 14980 17224 15008
rect 16982 14977 16994 14980
rect 16936 14971 16994 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 7834 14900 7840 14952
rect 7892 14940 7898 14952
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7892 14912 7941 14940
rect 7892 14900 7898 14912
rect 7929 14909 7941 14912
rect 7975 14940 7987 14943
rect 7975 14912 8432 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 6963 14844 7696 14872
rect 6963 14841 6975 14844
rect 6917 14835 6975 14841
rect 2685 14807 2743 14813
rect 2685 14773 2697 14807
rect 2731 14804 2743 14807
rect 2774 14804 2780 14816
rect 2731 14776 2780 14804
rect 2731 14773 2743 14776
rect 2685 14767 2743 14773
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 3326 14804 3332 14816
rect 3287 14776 3332 14804
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 4246 14804 4252 14816
rect 4207 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4488 14776 4629 14804
rect 4488 14764 4494 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 4617 14767 4675 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7248 14776 7297 14804
rect 7248 14764 7254 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 8404 14804 8432 14912
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16206 14940 16212 14952
rect 15528 14912 16212 14940
rect 15528 14900 15534 14912
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19536 14912 19901 14940
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 13446 14872 13452 14884
rect 10928 14844 13452 14872
rect 10928 14832 10934 14844
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 14384 14844 15884 14872
rect 10318 14804 10324 14816
rect 8404 14776 10324 14804
rect 7285 14767 7343 14773
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11054 14804 11060 14816
rect 10967 14776 11060 14804
rect 11054 14764 11060 14776
rect 11112 14804 11118 14816
rect 11238 14804 11244 14816
rect 11112 14776 11244 14804
rect 11112 14764 11118 14776
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11609 14807 11667 14813
rect 11609 14773 11621 14807
rect 11655 14804 11667 14807
rect 11698 14804 11704 14816
rect 11655 14776 11704 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 14384 14804 14412 14844
rect 13320 14776 14412 14804
rect 15197 14807 15255 14813
rect 13320 14764 13326 14776
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15243 14776 15669 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15657 14773 15669 14776
rect 15703 14804 15715 14807
rect 15746 14804 15752 14816
rect 15703 14776 15752 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 15856 14804 15884 14844
rect 19536 14816 19564 14912
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 16942 14804 16948 14816
rect 15856 14776 16948 14804
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 17368 14776 18061 14804
rect 17368 14764 17374 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18049 14767 18107 14773
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 18380 14776 18429 14804
rect 18380 14764 18386 14776
rect 18417 14773 18429 14776
rect 18463 14804 18475 14807
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18463 14776 18889 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 19518 14804 19524 14816
rect 19479 14776 19524 14804
rect 18877 14767 18935 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 20864 14776 21281 14804
rect 20864 14764 20870 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21269 14767 21327 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 5040 14572 5089 14600
rect 5040 14560 5046 14572
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 9766 14600 9772 14612
rect 5224 14572 9772 14600
rect 5224 14560 5230 14572
rect 9766 14560 9772 14572
rect 9824 14600 9830 14612
rect 10870 14600 10876 14612
rect 9824 14572 10876 14600
rect 9824 14560 9830 14572
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11885 14603 11943 14609
rect 11885 14600 11897 14603
rect 11020 14572 11897 14600
rect 11020 14560 11026 14572
rect 11885 14569 11897 14572
rect 11931 14569 11943 14603
rect 11885 14563 11943 14569
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13780 14572 14105 14600
rect 13780 14560 13786 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 15470 14600 15476 14612
rect 14093 14563 14151 14569
rect 14568 14572 15476 14600
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 3970 14532 3976 14544
rect 3844 14504 3976 14532
rect 3844 14492 3850 14504
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 9122 14532 9128 14544
rect 7024 14504 9128 14532
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14464 3479 14467
rect 3467 14436 4200 14464
rect 3467 14433 3479 14436
rect 3421 14427 3479 14433
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2777 14399 2835 14405
rect 2777 14396 2789 14399
rect 2179 14368 2789 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2777 14365 2789 14368
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3970 14396 3976 14408
rect 3099 14368 3976 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4172 14328 4200 14436
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 4304 14436 4353 14464
rect 4304 14424 4310 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5718 14464 5724 14476
rect 5132 14436 5724 14464
rect 5132 14424 5138 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 7024 14473 7052 14504
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 11974 14532 11980 14544
rect 11296 14504 11980 14532
rect 11296 14492 11302 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13446 14492 13452 14544
rect 13504 14532 13510 14544
rect 14568 14532 14596 14572
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15654 14560 15660 14612
rect 15712 14600 15718 14612
rect 16390 14600 16396 14612
rect 15712 14572 16396 14600
rect 15712 14560 15718 14572
rect 16390 14560 16396 14572
rect 16448 14600 16454 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 16448 14572 17141 14600
rect 16448 14560 16454 14572
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 17129 14563 17187 14569
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 18840 14572 19257 14600
rect 18840 14560 18846 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 19245 14563 19303 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 13504 14504 14596 14532
rect 13504 14492 13510 14504
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14433 7067 14467
rect 7190 14464 7196 14476
rect 7151 14436 7196 14464
rect 7009 14427 7067 14433
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9272 14436 10241 14464
rect 9272 14424 9278 14436
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8444 14368 8524 14396
rect 8444 14356 8450 14368
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 2792 14300 3832 14328
rect 4172 14300 4261 14328
rect 2792 14272 2820 14300
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2774 14220 2780 14272
rect 2832 14220 2838 14272
rect 3804 14269 3832 14300
rect 4249 14297 4261 14300
rect 4295 14328 4307 14331
rect 5166 14328 5172 14340
rect 4295 14300 5172 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 5445 14331 5503 14337
rect 5445 14297 5457 14331
rect 5491 14328 5503 14331
rect 5626 14328 5632 14340
rect 5491 14300 5632 14328
rect 5491 14297 5503 14300
rect 5445 14291 5503 14297
rect 5626 14288 5632 14300
rect 5684 14328 5690 14340
rect 6457 14331 6515 14337
rect 6457 14328 6469 14331
rect 5684 14300 6469 14328
rect 5684 14288 5690 14300
rect 6457 14297 6469 14300
rect 6503 14297 6515 14331
rect 6457 14291 6515 14297
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4157 14263 4215 14269
rect 4157 14260 4169 14263
rect 4120 14232 4169 14260
rect 4120 14220 4126 14232
rect 4157 14229 4169 14232
rect 4203 14260 4215 14263
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 4203 14232 5549 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 5537 14223 5595 14229
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5776 14232 6193 14260
rect 5776 14220 5782 14232
rect 6181 14229 6193 14232
rect 6227 14260 6239 14263
rect 6822 14260 6828 14272
rect 6227 14232 6828 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7653 14263 7711 14269
rect 7653 14229 7665 14263
rect 7699 14260 7711 14263
rect 8386 14260 8392 14272
rect 7699 14232 8392 14260
rect 7699 14229 7711 14232
rect 7653 14223 7711 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8496 14260 8524 14368
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 10134 14396 10140 14408
rect 8996 14368 10140 14396
rect 8996 14356 9002 14368
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 10502 14405 10508 14408
rect 10496 14396 10508 14405
rect 10463 14368 10508 14396
rect 10496 14359 10508 14368
rect 10502 14356 10508 14359
rect 10560 14356 10566 14408
rect 13265 14399 13323 14405
rect 10612 14368 13216 14396
rect 9306 14288 9312 14340
rect 9364 14328 9370 14340
rect 9490 14328 9496 14340
rect 9364 14300 9496 14328
rect 9364 14288 9370 14300
rect 9490 14288 9496 14300
rect 9548 14328 9554 14340
rect 10612 14328 10640 14368
rect 12998 14331 13056 14337
rect 12998 14328 13010 14331
rect 9548 14300 10640 14328
rect 10704 14300 13010 14328
rect 9548 14288 9554 14300
rect 8754 14260 8760 14272
rect 8496 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14260 8818 14272
rect 9950 14260 9956 14272
rect 8812 14232 9956 14260
rect 8812 14220 8818 14232
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10704 14260 10732 14300
rect 12998 14297 13010 14300
rect 13044 14297 13056 14331
rect 13188 14328 13216 14368
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 13538 14396 13544 14408
rect 13311 14368 13544 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15746 14396 15752 14408
rect 15519 14368 15752 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 16022 14405 16028 14408
rect 16016 14396 16028 14405
rect 15983 14368 16028 14396
rect 16016 14359 16028 14368
rect 16022 14356 16028 14359
rect 16080 14356 16086 14408
rect 18785 14399 18843 14405
rect 18785 14396 18797 14399
rect 18616 14368 18797 14396
rect 15206 14331 15264 14337
rect 15206 14328 15218 14331
rect 13188 14300 15218 14328
rect 12998 14291 13056 14297
rect 15206 14297 15218 14300
rect 15252 14297 15264 14331
rect 15206 14291 15264 14297
rect 15838 14288 15844 14340
rect 15896 14328 15902 14340
rect 18518 14331 18576 14337
rect 18518 14328 18530 14331
rect 15896 14300 18530 14328
rect 15896 14288 15902 14300
rect 18518 14297 18530 14300
rect 18564 14297 18576 14331
rect 18518 14291 18576 14297
rect 10100 14232 10732 14260
rect 11609 14263 11667 14269
rect 10100 14220 10106 14232
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 11790 14260 11796 14272
rect 11655 14232 11796 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 13538 14260 13544 14272
rect 12952 14232 13544 14260
rect 12952 14220 12958 14232
rect 13538 14220 13544 14232
rect 13596 14260 13602 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13596 14232 13645 14260
rect 13596 14220 13602 14232
rect 13633 14229 13645 14232
rect 13679 14260 13691 14263
rect 14458 14260 14464 14272
rect 13679 14232 14464 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 18322 14220 18328 14272
rect 18380 14260 18386 14272
rect 18616 14260 18644 14368
rect 18785 14365 18797 14368
rect 18831 14396 18843 14399
rect 19334 14396 19340 14408
rect 18831 14368 19340 14396
rect 18831 14365 18843 14368
rect 18785 14359 18843 14365
rect 19334 14356 19340 14368
rect 19392 14396 19398 14408
rect 19518 14396 19524 14408
rect 19392 14368 19524 14396
rect 19392 14356 19398 14368
rect 19518 14356 19524 14368
rect 19576 14396 19582 14408
rect 20622 14396 20628 14408
rect 19576 14368 20628 14396
rect 19576 14356 19582 14368
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20772 14368 20913 14396
rect 20772 14356 20778 14368
rect 20901 14365 20913 14368
rect 20947 14396 20959 14399
rect 21266 14396 21272 14408
rect 20947 14368 21272 14396
rect 20947 14365 20959 14368
rect 20901 14359 20959 14365
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 19978 14288 19984 14340
rect 20036 14328 20042 14340
rect 20346 14328 20352 14340
rect 20404 14337 20410 14340
rect 20036 14300 20352 14328
rect 20036 14288 20042 14300
rect 20346 14288 20352 14300
rect 20404 14328 20416 14337
rect 20404 14300 20449 14328
rect 20404 14291 20416 14300
rect 20404 14288 20410 14291
rect 18380 14232 18644 14260
rect 18380 14220 18386 14232
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4430 14056 4436 14068
rect 4391 14028 4436 14056
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 5316 14028 5549 14056
rect 5316 14016 5322 14028
rect 5537 14025 5549 14028
rect 5583 14056 5595 14059
rect 5583 14028 12434 14056
rect 5583 14025 5595 14028
rect 5537 14019 5595 14025
rect 3697 13991 3755 13997
rect 3697 13957 3709 13991
rect 3743 13988 3755 13991
rect 4062 13988 4068 14000
rect 3743 13960 4068 13988
rect 3743 13957 3755 13960
rect 3697 13951 3755 13957
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 4338 13988 4344 14000
rect 4299 13960 4344 13988
rect 4338 13948 4344 13960
rect 4396 13948 4402 14000
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 6917 13991 6975 13997
rect 6917 13988 6929 13991
rect 5868 13960 6929 13988
rect 5868 13948 5874 13960
rect 6917 13957 6929 13960
rect 6963 13988 6975 13991
rect 8113 13991 8171 13997
rect 8113 13988 8125 13991
rect 6963 13960 8125 13988
rect 6963 13957 6975 13960
rect 6917 13951 6975 13957
rect 8113 13957 8125 13960
rect 8159 13988 8171 13991
rect 8754 13988 8760 14000
rect 8159 13960 8760 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 12406 13988 12434 14028
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 12860 14028 14289 14056
rect 12860 14016 12866 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 14292 13988 14320 14019
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15344 14028 15945 14056
rect 15344 14016 15350 14028
rect 15933 14025 15945 14028
rect 15979 14056 15991 14059
rect 16022 14056 16028 14068
rect 15979 14028 16028 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 18966 14056 18972 14068
rect 18927 14028 18972 14056
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19334 14056 19340 14068
rect 19295 14028 19340 14056
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19760 14028 19901 14056
rect 19760 14016 19766 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 19889 14019 19947 14025
rect 14798 13991 14856 13997
rect 14798 13988 14810 13991
rect 9232 13960 11008 13988
rect 12406 13960 13308 13988
rect 14292 13960 14810 13988
rect 9232 13932 9260 13960
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2409 13923 2467 13929
rect 2409 13920 2421 13923
rect 1995 13892 2421 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2409 13889 2421 13892
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 2590 13880 2596 13932
rect 2648 13920 2654 13932
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2648 13892 2697 13920
rect 2648 13880 2654 13892
rect 2685 13889 2697 13892
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 3844 13892 6837 13920
rect 3844 13880 3850 13892
rect 6825 13889 6837 13892
rect 6871 13920 6883 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 6871 13892 8401 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 8389 13889 8401 13892
rect 8435 13920 8447 13923
rect 8938 13920 8944 13932
rect 8435 13892 8944 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9490 13929 9496 13932
rect 9484 13920 9496 13929
rect 9451 13892 9496 13920
rect 9484 13883 9496 13892
rect 9490 13880 9496 13883
rect 9548 13880 9554 13932
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10100 13892 10272 13920
rect 10100 13880 10106 13892
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5074 13852 5080 13864
rect 4663 13824 5080 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5810 13852 5816 13864
rect 5771 13824 5816 13852
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7147 13824 7757 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 10244 13852 10272 13892
rect 10980 13861 11008 13960
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 13153 13923 13211 13929
rect 13153 13920 13165 13923
rect 11848 13892 13165 13920
rect 11848 13880 11854 13892
rect 13153 13889 13165 13892
rect 13199 13889 13211 13923
rect 13280 13920 13308 13960
rect 14798 13957 14810 13960
rect 14844 13957 14856 13991
rect 14798 13951 14856 13957
rect 17856 13991 17914 13997
rect 17856 13957 17868 13991
rect 17902 13988 17914 13991
rect 19720 13988 19748 14016
rect 17902 13960 19748 13988
rect 17902 13957 17914 13960
rect 17856 13951 17914 13957
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20680 13960 21312 13988
rect 20680 13948 20686 13960
rect 17218 13920 17224 13932
rect 13280 13892 17224 13920
rect 13153 13883 13211 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 17586 13920 17592 13932
rect 17359 13892 17592 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 10965 13855 11023 13861
rect 10244 13824 10640 13852
rect 7745 13815 7803 13821
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 7466 13784 7472 13796
rect 4120 13756 7472 13784
rect 4120 13744 4126 13756
rect 7466 13744 7472 13756
rect 7524 13744 7530 13796
rect 7760 13784 7788 13815
rect 10612 13793 10640 13824
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11698 13852 11704 13864
rect 11011 13824 11704 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11698 13812 11704 13824
rect 11756 13852 11762 13864
rect 12894 13852 12900 13864
rect 11756 13824 12900 13852
rect 11756 13812 11762 13824
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 10597 13787 10655 13793
rect 7760 13756 9260 13784
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 5074 13716 5080 13728
rect 5035 13688 5080 13716
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 5718 13676 5724 13728
rect 5776 13716 5782 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 5776 13688 6469 13716
rect 5776 13676 5782 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 9232 13716 9260 13756
rect 10597 13753 10609 13787
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 10134 13716 10140 13728
rect 9232 13688 10140 13716
rect 6457 13679 6515 13685
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 14458 13676 14464 13728
rect 14516 13716 14522 13728
rect 14568 13716 14596 13815
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16022 13852 16028 13864
rect 15804 13824 16028 13852
rect 15804 13812 15810 13824
rect 16022 13812 16028 13824
rect 16080 13852 16086 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16080 13824 16313 13852
rect 16080 13812 16086 13824
rect 16301 13821 16313 13824
rect 16347 13852 16359 13855
rect 17328 13852 17356 13883
rect 17586 13880 17592 13892
rect 17644 13920 17650 13932
rect 18322 13920 18328 13932
rect 17644 13892 18328 13920
rect 17644 13880 17650 13892
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 19702 13880 19708 13932
rect 19760 13920 19766 13932
rect 20990 13920 20996 13932
rect 21048 13929 21054 13932
rect 21284 13929 21312 13960
rect 19760 13892 20996 13920
rect 19760 13880 19766 13892
rect 20990 13880 20996 13892
rect 21048 13920 21060 13929
rect 21269 13923 21327 13929
rect 21048 13892 21093 13920
rect 21048 13883 21060 13892
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21048 13880 21054 13883
rect 16347 13824 17356 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 15764 13716 15792 13812
rect 14516 13688 15792 13716
rect 14516 13676 14522 13688
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 1854 13512 1860 13524
rect 1719 13484 1860 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3476 13484 3801 13512
rect 3476 13472 3482 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6052 13484 6469 13512
rect 6052 13472 6058 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 6457 13475 6515 13481
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8168 13484 10364 13512
rect 8168 13472 8174 13484
rect 6181 13447 6239 13453
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 6546 13444 6552 13456
rect 6227 13416 6552 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 10336 13444 10364 13484
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10560 13484 10793 13512
rect 10560 13472 10566 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 14458 13512 14464 13524
rect 14419 13484 14464 13512
rect 10781 13475 10839 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17092 13484 17417 13512
rect 17092 13472 17098 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 17644 13484 17693 13512
rect 17644 13472 17650 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 21082 13512 21088 13524
rect 21043 13484 21088 13512
rect 17681 13475 17739 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 14550 13444 14556 13456
rect 6932 13416 8156 13444
rect 10336 13416 14556 13444
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 4430 13376 4436 13388
rect 4391 13348 4436 13376
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 6932 13376 6960 13416
rect 5675 13348 6960 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 7006 13336 7012 13388
rect 7064 13376 7070 13388
rect 8128 13385 8156 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 8113 13379 8171 13385
rect 7064 13348 7109 13376
rect 7064 13336 7070 13348
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8159 13348 9076 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 5810 13308 5816 13320
rect 5771 13280 5816 13308
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6880 13280 6929 13308
rect 6880 13268 6886 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 2746 13212 4169 13240
rect 2038 13172 2044 13184
rect 1999 13144 2044 13172
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2188 13144 2233 13172
rect 2188 13132 2194 13144
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2746 13172 2774 13212
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 5169 13243 5227 13249
rect 5169 13240 5181 13243
rect 4157 13203 4215 13209
rect 4448 13212 5181 13240
rect 4448 13184 4476 13212
rect 5169 13209 5181 13212
rect 5215 13240 5227 13243
rect 5442 13240 5448 13252
rect 5215 13212 5448 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 5442 13200 5448 13212
rect 5500 13240 5506 13252
rect 5721 13243 5779 13249
rect 5721 13240 5733 13243
rect 5500 13212 5733 13240
rect 5500 13200 5506 13212
rect 5721 13209 5733 13212
rect 5767 13209 5779 13243
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 5721 13203 5779 13209
rect 5828 13212 6868 13240
rect 5828 13184 5856 13212
rect 4246 13172 4252 13184
rect 2556 13144 2774 13172
rect 4207 13144 4252 13172
rect 2556 13132 2562 13144
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4430 13132 4436 13184
rect 4488 13132 4494 13184
rect 5810 13132 5816 13184
rect 5868 13132 5874 13184
rect 6840 13181 6868 13212
rect 7852 13212 8953 13240
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13141 6883 13175
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 6825 13135 6883 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7852 13181 7880 13212
rect 8941 13209 8953 13212
rect 8987 13209 8999 13243
rect 8941 13203 8999 13209
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7800 13144 7849 13172
rect 7800 13132 7806 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 7929 13175 7987 13181
rect 7929 13141 7941 13175
rect 7975 13172 7987 13175
rect 8110 13172 8116 13184
rect 7975 13144 8116 13172
rect 7975 13141 7987 13144
rect 7929 13135 7987 13141
rect 8110 13132 8116 13144
rect 8168 13172 8174 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8168 13144 8493 13172
rect 8168 13132 8174 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 9048 13172 9076 13348
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9272 13348 9413 13376
rect 9272 13336 9278 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 12406 13348 16160 13376
rect 12406 13308 12434 13348
rect 16022 13308 16028 13320
rect 9232 13280 12434 13308
rect 15983 13280 16028 13308
rect 9232 13252 9260 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16132 13308 16160 13348
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 16132 13280 18797 13308
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 18785 13271 18843 13277
rect 20180 13280 20637 13308
rect 9214 13200 9220 13252
rect 9272 13200 9278 13252
rect 9668 13243 9726 13249
rect 9668 13209 9680 13243
rect 9714 13240 9726 13243
rect 9858 13240 9864 13252
rect 9714 13212 9864 13240
rect 9714 13209 9726 13212
rect 9668 13203 9726 13209
rect 9858 13200 9864 13212
rect 9916 13240 9922 13252
rect 12250 13240 12256 13252
rect 9916 13212 12256 13240
rect 9916 13200 9922 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 16292 13243 16350 13249
rect 16292 13209 16304 13243
rect 16338 13240 16350 13243
rect 16390 13240 16396 13252
rect 16338 13212 16396 13240
rect 16338 13209 16350 13212
rect 16292 13203 16350 13209
rect 16390 13200 16396 13212
rect 16448 13200 16454 13252
rect 18800 13240 18828 13271
rect 20180 13252 20208 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 18800 13212 20116 13240
rect 10042 13172 10048 13184
rect 9048 13144 10048 13172
rect 8481 13135 8539 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 11149 13175 11207 13181
rect 11149 13141 11161 13175
rect 11195 13172 11207 13175
rect 11698 13172 11704 13184
rect 11195 13144 11704 13172
rect 11195 13141 11207 13144
rect 11149 13135 11207 13141
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 17126 13132 17132 13184
rect 17184 13172 17190 13184
rect 17310 13172 17316 13184
rect 17184 13144 17316 13172
rect 17184 13132 17190 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 18196 13144 19257 13172
rect 18196 13132 18202 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 20088 13172 20116 13212
rect 20162 13200 20168 13252
rect 20220 13200 20226 13252
rect 20380 13243 20438 13249
rect 20380 13209 20392 13243
rect 20426 13240 20438 13243
rect 20806 13240 20812 13252
rect 20426 13212 20812 13240
rect 20426 13209 20438 13212
rect 20380 13203 20438 13209
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 20916 13172 20944 13271
rect 20088 13144 20944 13172
rect 19245 13135 19303 13141
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 2096 12940 2421 12968
rect 2096 12928 2102 12940
rect 2409 12937 2421 12940
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4304 12940 5273 12968
rect 4304 12928 4310 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5261 12931 5319 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6730 12968 6736 12980
rect 6236 12940 6736 12968
rect 6236 12928 6242 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7432 12940 7665 12968
rect 7432 12928 7438 12940
rect 7653 12937 7665 12940
rect 7699 12968 7711 12971
rect 8570 12968 8576 12980
rect 7699 12940 8576 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 8570 12928 8576 12940
rect 8628 12968 8634 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8628 12940 8677 12968
rect 8628 12928 8634 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 8665 12931 8723 12937
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9306 12968 9312 12980
rect 9263 12940 9312 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10410 12968 10416 12980
rect 10008 12940 10416 12968
rect 10008 12928 10014 12940
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10928 12940 10977 12968
rect 10928 12928 10934 12940
rect 10965 12937 10977 12940
rect 11011 12968 11023 12971
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11011 12940 11621 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 11609 12937 11621 12940
rect 11655 12968 11667 12971
rect 11698 12968 11704 12980
rect 11655 12940 11704 12968
rect 11655 12937 11667 12940
rect 11609 12931 11667 12937
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 13906 12968 13912 12980
rect 12406 12940 13912 12968
rect 4338 12860 4344 12912
rect 4396 12900 4402 12912
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4396 12872 4537 12900
rect 4396 12860 4402 12872
rect 4525 12869 4537 12872
rect 4571 12869 4583 12903
rect 4525 12863 4583 12869
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 8110 12900 8116 12912
rect 4856 12872 8116 12900
rect 4856 12860 4862 12872
rect 8110 12860 8116 12872
rect 8168 12900 8174 12912
rect 8297 12903 8355 12909
rect 8297 12900 8309 12903
rect 8168 12872 8309 12900
rect 8168 12860 8174 12872
rect 8297 12869 8309 12872
rect 8343 12869 8355 12903
rect 8297 12863 8355 12869
rect 10226 12860 10232 12912
rect 10284 12900 10290 12912
rect 10330 12903 10388 12909
rect 10330 12900 10342 12903
rect 10284 12872 10342 12900
rect 10284 12860 10290 12872
rect 10330 12869 10342 12872
rect 10376 12869 10388 12903
rect 12406 12900 12434 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12937 14151 12971
rect 14093 12931 14151 12937
rect 15841 12971 15899 12977
rect 15841 12937 15853 12971
rect 15887 12968 15899 12971
rect 16022 12968 16028 12980
rect 15887 12940 16028 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 14108 12900 14136 12931
rect 10330 12863 10388 12869
rect 11072 12872 12434 12900
rect 12912 12872 14136 12900
rect 15228 12903 15286 12909
rect 1670 12792 1676 12844
rect 1728 12832 1734 12844
rect 2041 12835 2099 12841
rect 2041 12832 2053 12835
rect 1728 12804 2053 12832
rect 1728 12792 1734 12804
rect 2041 12801 2053 12804
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 2740 12804 3709 12832
rect 2740 12792 2746 12804
rect 3697 12801 3709 12804
rect 3743 12832 3755 12835
rect 4982 12832 4988 12844
rect 3743 12804 4988 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 1946 12764 1952 12776
rect 1907 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4614 12764 4620 12776
rect 3651 12736 4620 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 3528 12696 3556 12727
rect 4614 12724 4620 12736
rect 4672 12764 4678 12776
rect 4798 12764 4804 12776
rect 4672 12736 4804 12764
rect 4672 12724 4678 12736
rect 4798 12724 4804 12736
rect 4856 12764 4862 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4856 12736 4905 12764
rect 4856 12724 4862 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 5644 12708 5672 12795
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 7006 12832 7012 12844
rect 6144 12804 7012 12832
rect 6144 12792 6150 12804
rect 7006 12792 7012 12804
rect 7064 12832 7070 12844
rect 10597 12835 10655 12841
rect 7064 12804 10548 12832
rect 7064 12792 7070 12804
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 5994 12764 6000 12776
rect 5951 12736 6000 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 7742 12764 7748 12776
rect 6564 12736 7748 12764
rect 3970 12696 3976 12708
rect 3528 12668 3976 12696
rect 3970 12656 3976 12668
rect 4028 12696 4034 12708
rect 4338 12696 4344 12708
rect 4028 12668 4344 12696
rect 4028 12656 4034 12668
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 5626 12656 5632 12708
rect 5684 12656 5690 12708
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4246 12628 4252 12640
rect 4111 12600 4252 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 5258 12588 5264 12640
rect 5316 12628 5322 12640
rect 6564 12637 6592 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 10520 12764 10548 12804
rect 10597 12801 10609 12835
rect 10643 12832 10655 12835
rect 10870 12832 10876 12844
rect 10643 12804 10876 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11072 12764 11100 12872
rect 12912 12832 12940 12872
rect 15228 12869 15240 12903
rect 15274 12900 15286 12903
rect 15654 12900 15660 12912
rect 15274 12872 15660 12900
rect 15274 12869 15286 12872
rect 15228 12863 15286 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 10520 12736 11100 12764
rect 12406 12804 12940 12832
rect 13561 12835 13619 12841
rect 7837 12727 7895 12733
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7852 12696 7880 12727
rect 12406 12696 12434 12804
rect 13561 12801 13573 12835
rect 13607 12832 13619 12835
rect 14458 12832 14464 12844
rect 13607 12804 14464 12832
rect 13607 12801 13619 12804
rect 13561 12795 13619 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 15746 12832 15752 12844
rect 15519 12804 15752 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15746 12792 15752 12804
rect 15804 12832 15810 12844
rect 15856 12832 15884 12931
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 19058 12928 19064 12980
rect 19116 12968 19122 12980
rect 19245 12971 19303 12977
rect 19245 12968 19257 12971
rect 19116 12940 19257 12968
rect 19116 12928 19122 12940
rect 19245 12937 19257 12940
rect 19291 12937 19303 12971
rect 19245 12931 19303 12937
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19576 12940 20085 12968
rect 19576 12928 19582 12940
rect 20073 12937 20085 12940
rect 20119 12968 20131 12971
rect 20162 12968 20168 12980
rect 20119 12940 20168 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20254 12928 20260 12980
rect 20312 12968 20318 12980
rect 20533 12971 20591 12977
rect 20533 12968 20545 12971
rect 20312 12940 20545 12968
rect 20312 12928 20318 12940
rect 20533 12937 20545 12940
rect 20579 12937 20591 12971
rect 20533 12931 20591 12937
rect 19702 12900 19708 12912
rect 19663 12872 19708 12900
rect 19702 12860 19708 12872
rect 19760 12900 19766 12912
rect 19760 12872 20300 12900
rect 19760 12860 19766 12872
rect 20272 12844 20300 12872
rect 15804 12804 15884 12832
rect 15804 12792 15810 12804
rect 17586 12792 17592 12844
rect 17644 12832 17650 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17644 12804 17877 12832
rect 17644 12792 17650 12804
rect 17865 12801 17877 12804
rect 17911 12801 17923 12835
rect 17865 12795 17923 12801
rect 18132 12835 18190 12841
rect 18132 12801 18144 12835
rect 18178 12832 18190 12835
rect 19794 12832 19800 12844
rect 18178 12804 19800 12832
rect 18178 12801 18190 12804
rect 18132 12795 18190 12801
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 20254 12792 20260 12844
rect 20312 12792 20318 12844
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12832 20959 12835
rect 21266 12832 21272 12844
rect 20947 12804 21272 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 13814 12764 13820 12776
rect 13775 12736 13820 12764
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 20990 12764 20996 12776
rect 20951 12736 20996 12764
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21085 12767 21143 12773
rect 21085 12733 21097 12767
rect 21131 12733 21143 12767
rect 21085 12727 21143 12733
rect 6788 12668 7880 12696
rect 10612 12668 12434 12696
rect 6788 12656 6794 12668
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 5316 12600 6561 12628
rect 5316 12588 5322 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 6549 12591 6607 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 8202 12588 8208 12640
rect 8260 12628 8266 12640
rect 9306 12628 9312 12640
rect 8260 12600 9312 12628
rect 8260 12588 8266 12600
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10612 12628 10640 12668
rect 19978 12656 19984 12708
rect 20036 12696 20042 12708
rect 21100 12696 21128 12727
rect 20036 12668 21128 12696
rect 20036 12656 20042 12668
rect 12434 12628 12440 12640
rect 10284 12600 10640 12628
rect 12395 12600 12440 12628
rect 10284 12588 10290 12600
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 15286 12628 15292 12640
rect 13964 12600 15292 12628
rect 13964 12588 13970 12600
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4154 12424 4160 12436
rect 3927 12396 4160 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5902 12424 5908 12436
rect 5684 12396 5908 12424
rect 5684 12384 5690 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6880 12396 6929 12424
rect 6880 12384 6886 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 11790 12424 11796 12436
rect 6917 12387 6975 12393
rect 7024 12396 11796 12424
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 7024 12356 7052 12396
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 12250 12424 12256 12436
rect 12211 12396 12256 12424
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 14458 12424 14464 12436
rect 14419 12396 14464 12424
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 17405 12427 17463 12433
rect 17405 12393 17417 12427
rect 17451 12424 17463 12427
rect 17586 12424 17592 12436
rect 17451 12396 17592 12424
rect 17451 12393 17463 12396
rect 17405 12387 17463 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20346 12424 20352 12436
rect 20119 12396 20352 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21269 12427 21327 12433
rect 21269 12424 21281 12427
rect 21048 12396 21281 12424
rect 21048 12384 21054 12396
rect 21269 12393 21281 12396
rect 21315 12393 21327 12427
rect 21269 12387 21327 12393
rect 8662 12356 8668 12368
rect 3108 12328 7052 12356
rect 7392 12328 8668 12356
rect 3108 12316 3114 12328
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 2682 12288 2688 12300
rect 2547 12260 2688 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4120 12260 4445 12288
rect 4120 12248 4126 12260
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6822 12288 6828 12300
rect 6135 12260 6828 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6822 12248 6828 12260
rect 6880 12288 6886 12300
rect 7392 12288 7420 12328
rect 8662 12316 8668 12328
rect 8720 12316 8726 12368
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 9217 12359 9275 12365
rect 9217 12356 9229 12359
rect 9180 12328 9229 12356
rect 9180 12316 9186 12328
rect 9217 12325 9229 12328
rect 9263 12325 9275 12359
rect 9217 12319 9275 12325
rect 7558 12288 7564 12300
rect 6880 12260 7420 12288
rect 7519 12260 7564 12288
rect 6880 12248 6886 12260
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2774 12220 2780 12232
rect 2363 12192 2780 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2774 12180 2780 12192
rect 2832 12180 2838 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6178 12220 6184 12232
rect 5960 12192 6184 12220
rect 5960 12180 5966 12192
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 8110 12220 8116 12232
rect 7331 12192 8116 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 9232 12220 9260 12319
rect 13170 12316 13176 12368
rect 13228 12356 13234 12368
rect 15654 12356 15660 12368
rect 13228 12328 15660 12356
rect 13228 12316 13234 12328
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 10597 12291 10655 12297
rect 10597 12257 10609 12291
rect 10643 12288 10655 12291
rect 10870 12288 10876 12300
rect 10643 12260 10876 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 20806 12288 20812 12300
rect 20763 12260 20812 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 12621 12223 12679 12229
rect 9232 12192 10548 12220
rect 1762 12112 1768 12164
rect 1820 12152 1826 12164
rect 1820 12124 9352 12152
rect 1820 12112 1826 12124
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 1857 12087 1915 12093
rect 1857 12053 1869 12087
rect 1903 12084 1915 12087
rect 2038 12084 2044 12096
rect 1903 12056 2044 12084
rect 1903 12053 1915 12056
rect 1857 12047 1915 12053
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 2869 12087 2927 12093
rect 2869 12084 2881 12087
rect 2740 12056 2881 12084
rect 2740 12044 2746 12056
rect 2869 12053 2881 12056
rect 2915 12053 2927 12087
rect 3234 12084 3240 12096
rect 3195 12056 3240 12084
rect 2869 12047 2927 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 3568 12056 4261 12084
rect 3568 12044 3574 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4890 12084 4896 12096
rect 4396 12056 4441 12084
rect 4851 12056 4896 12084
rect 4396 12044 4402 12056
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5258 12084 5264 12096
rect 5219 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6914 12084 6920 12096
rect 6595 12056 6920 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 7156 12056 7389 12084
rect 7156 12044 7162 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 7616 12056 8125 12084
rect 7616 12044 7622 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 8260 12056 8493 12084
rect 8260 12044 8266 12056
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 9324 12084 9352 12124
rect 10318 12112 10324 12164
rect 10376 12161 10382 12164
rect 10376 12152 10388 12161
rect 10520 12152 10548 12192
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 13814 12220 13820 12232
rect 12667 12192 13820 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 13814 12180 13820 12192
rect 13872 12220 13878 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13872 12192 14197 12220
rect 13872 12180 13878 12192
rect 14185 12189 14197 12192
rect 14231 12220 14243 12223
rect 14918 12220 14924 12232
rect 14231 12192 14924 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14918 12180 14924 12192
rect 14976 12220 14982 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 14976 12192 15669 12220
rect 14976 12180 14982 12192
rect 15657 12189 15669 12192
rect 15703 12220 15715 12223
rect 15746 12220 15752 12232
rect 15703 12192 15752 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 20254 12220 20260 12232
rect 20215 12192 20260 12220
rect 20254 12180 20260 12192
rect 20312 12180 20318 12232
rect 11118 12155 11176 12161
rect 11118 12152 11130 12155
rect 10376 12124 10421 12152
rect 10520 12124 11130 12152
rect 10376 12115 10388 12124
rect 11118 12121 11130 12124
rect 11164 12121 11176 12155
rect 13262 12152 13268 12164
rect 11118 12115 11176 12121
rect 12406 12124 13268 12152
rect 10376 12112 10382 12115
rect 12406 12084 12434 12124
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 15286 12112 15292 12164
rect 15344 12152 15350 12164
rect 15924 12155 15982 12161
rect 15924 12152 15936 12155
rect 15344 12124 15936 12152
rect 15344 12112 15350 12124
rect 15924 12121 15936 12124
rect 15970 12152 15982 12155
rect 17586 12152 17592 12164
rect 15970 12124 17592 12152
rect 15970 12121 15982 12124
rect 15924 12115 15982 12121
rect 17586 12112 17592 12124
rect 17644 12152 17650 12164
rect 17681 12155 17739 12161
rect 17681 12152 17693 12155
rect 17644 12124 17693 12152
rect 17644 12112 17650 12124
rect 17681 12121 17693 12124
rect 17727 12121 17739 12155
rect 17681 12115 17739 12121
rect 19337 12155 19395 12161
rect 19337 12121 19349 12155
rect 19383 12152 19395 12155
rect 19702 12152 19708 12164
rect 19383 12124 19708 12152
rect 19383 12121 19395 12124
rect 19337 12115 19395 12121
rect 19702 12112 19708 12124
rect 19760 12152 19766 12164
rect 19886 12152 19892 12164
rect 19760 12124 19892 12152
rect 19760 12112 19766 12124
rect 19886 12112 19892 12124
rect 19944 12152 19950 12164
rect 20809 12155 20867 12161
rect 20809 12152 20821 12155
rect 19944 12124 20821 12152
rect 19944 12112 19950 12124
rect 20809 12121 20821 12124
rect 20855 12121 20867 12155
rect 20809 12115 20867 12121
rect 9324 12056 12434 12084
rect 8481 12047 8539 12053
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 17000 12056 17049 12084
rect 17000 12044 17006 12056
rect 17037 12053 17049 12056
rect 17083 12084 17095 12087
rect 17218 12084 17224 12096
rect 17083 12056 17224 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18506 12084 18512 12096
rect 18196 12056 18512 12084
rect 18196 12044 18202 12056
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19610 12084 19616 12096
rect 19571 12056 19616 12084
rect 19610 12044 19616 12056
rect 19668 12084 19674 12096
rect 19978 12084 19984 12096
rect 19668 12056 19984 12084
rect 19668 12044 19674 12056
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 20990 12084 20996 12096
rect 20947 12056 20996 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2188 11852 2421 11880
rect 2188 11840 2194 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3234 11880 3240 11892
rect 3099 11852 3240 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 3510 11880 3516 11892
rect 3471 11852 3516 11880
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4246 11880 4252 11892
rect 4207 11852 4252 11880
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4396 11852 5273 11880
rect 4396 11840 4402 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 6638 11840 6644 11892
rect 6696 11880 6702 11892
rect 7098 11880 7104 11892
rect 6696 11852 7104 11880
rect 6696 11840 6702 11852
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 7466 11880 7472 11892
rect 7239 11852 7472 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 9490 11880 9496 11892
rect 7708 11852 9496 11880
rect 7708 11840 7714 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 11698 11880 11704 11892
rect 9600 11852 11704 11880
rect 1854 11772 1860 11824
rect 1912 11812 1918 11824
rect 4893 11815 4951 11821
rect 4893 11812 4905 11815
rect 1912 11784 4905 11812
rect 1912 11772 1918 11784
rect 4893 11781 4905 11784
rect 4939 11812 4951 11815
rect 5629 11815 5687 11821
rect 5629 11812 5641 11815
rect 4939 11784 5641 11812
rect 4939 11781 4951 11784
rect 4893 11775 4951 11781
rect 5629 11781 5641 11784
rect 5675 11812 5687 11815
rect 5718 11812 5724 11824
rect 5675 11784 5724 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 5718 11772 5724 11784
rect 5776 11772 5782 11824
rect 6546 11772 6552 11824
rect 6604 11812 6610 11824
rect 7285 11815 7343 11821
rect 7285 11812 7297 11815
rect 6604 11784 7297 11812
rect 6604 11772 6610 11784
rect 7285 11781 7297 11784
rect 7331 11781 7343 11815
rect 7285 11775 7343 11781
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 8202 11812 8208 11824
rect 7984 11784 8208 11812
rect 7984 11772 7990 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 8662 11812 8668 11824
rect 8575 11784 8668 11812
rect 8662 11772 8668 11784
rect 8720 11812 8726 11824
rect 9600 11812 9628 11852
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 13170 11880 13176 11892
rect 11808 11852 12204 11880
rect 13131 11852 13176 11880
rect 11146 11812 11152 11824
rect 8720 11784 9628 11812
rect 10060 11784 11152 11812
rect 8720 11772 8726 11784
rect 3142 11744 3148 11756
rect 3103 11716 3148 11744
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4982 11744 4988 11756
rect 4203 11716 4988 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 6822 11744 6828 11756
rect 5736 11716 6828 11744
rect 1762 11676 1768 11688
rect 1723 11648 1768 11676
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 1949 11639 2007 11645
rect 1964 11608 1992 11639
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11676 4491 11679
rect 5258 11676 5264 11688
rect 4479 11648 5264 11676
rect 4479 11645 4491 11648
rect 4433 11639 4491 11645
rect 3789 11611 3847 11617
rect 3789 11608 3801 11611
rect 1964 11580 3801 11608
rect 3789 11577 3801 11580
rect 3835 11577 3847 11611
rect 3789 11571 3847 11577
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2682 11540 2688 11552
rect 2188 11512 2688 11540
rect 2188 11500 2194 11512
rect 2682 11500 2688 11512
rect 2740 11540 2746 11552
rect 4448 11540 4476 11639
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5736 11685 5764 11716
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 10060 11744 10088 11784
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11808 11812 11836 11852
rect 11664 11784 11836 11812
rect 11664 11772 11670 11784
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 12038 11815 12096 11821
rect 12038 11812 12050 11815
rect 11940 11784 12050 11812
rect 11940 11772 11946 11784
rect 12038 11781 12050 11784
rect 12084 11781 12096 11815
rect 12176 11812 12204 11852
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13280 11852 15332 11880
rect 13280 11812 13308 11852
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 12176 11784 13308 11812
rect 13372 11784 13553 11812
rect 12038 11775 12096 11781
rect 7116 11716 10088 11744
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 6086 11676 6092 11688
rect 5951 11648 6092 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 5626 11568 5632 11620
rect 5684 11608 5690 11620
rect 5920 11608 5948 11639
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 7116 11685 7144 11716
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10606 11747 10664 11753
rect 10606 11744 10618 11747
rect 10192 11716 10618 11744
rect 10192 11704 10198 11716
rect 10606 11713 10618 11716
rect 10652 11713 10664 11747
rect 10870 11744 10876 11756
rect 10831 11716 10876 11744
rect 10606 11707 10664 11713
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 13372 11744 13400 11784
rect 13541 11781 13553 11784
rect 13587 11812 13599 11815
rect 13814 11812 13820 11824
rect 13587 11784 13820 11812
rect 13587 11781 13599 11784
rect 13541 11775 13599 11781
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 15166 11815 15224 11821
rect 15166 11812 15178 11815
rect 14884 11784 15178 11812
rect 14884 11772 14890 11784
rect 15166 11781 15178 11784
rect 15212 11781 15224 11815
rect 15304 11812 15332 11852
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 18598 11880 18604 11892
rect 16356 11852 18604 11880
rect 16356 11840 16362 11852
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 20162 11880 20168 11892
rect 19751 11852 20168 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 20162 11840 20168 11852
rect 20220 11880 20226 11892
rect 20622 11880 20628 11892
rect 20220 11852 20628 11880
rect 20220 11840 20226 11852
rect 20622 11840 20628 11852
rect 20680 11880 20686 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 20680 11852 21189 11880
rect 20680 11840 20686 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 18224 11815 18282 11821
rect 15304 11784 18175 11812
rect 15166 11775 15224 11781
rect 11839 11716 13400 11744
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 18046 11744 18052 11756
rect 13504 11716 18052 11744
rect 13504 11704 13510 11716
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18147 11744 18175 11784
rect 18224 11781 18236 11815
rect 18270 11812 18282 11815
rect 19058 11812 19064 11824
rect 18270 11784 19064 11812
rect 18270 11781 18282 11784
rect 18224 11775 18282 11781
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 20254 11772 20260 11824
rect 20312 11812 20318 11824
rect 20717 11815 20775 11821
rect 20717 11812 20729 11815
rect 20312 11784 20729 11812
rect 20312 11772 20318 11784
rect 20717 11781 20729 11784
rect 20763 11781 20775 11815
rect 20717 11775 20775 11781
rect 20438 11744 20444 11756
rect 18147 11716 19334 11744
rect 20399 11716 20444 11744
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7926 11676 7932 11688
rect 7887 11648 7932 11676
rect 7101 11639 7159 11645
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 17957 11679 18015 11685
rect 17957 11676 17969 11679
rect 17920 11648 17969 11676
rect 17920 11636 17926 11648
rect 17957 11645 17969 11648
rect 18003 11645 18015 11679
rect 19306 11676 19334 11716
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20714 11676 20720 11688
rect 19306 11648 20720 11676
rect 17957 11639 18015 11645
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 11606 11608 11612 11620
rect 5684 11580 5948 11608
rect 6012 11580 8524 11608
rect 5684 11568 5690 11580
rect 2740 11512 4476 11540
rect 2740 11500 2746 11512
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 6012 11540 6040 11580
rect 8496 11552 8524 11580
rect 10888 11580 11612 11608
rect 4672 11512 6040 11540
rect 4672 11500 4678 11512
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 6144 11512 6469 11540
rect 6144 11500 6150 11512
rect 6457 11509 6469 11512
rect 6503 11540 6515 11543
rect 6546 11540 6552 11552
rect 6503 11512 6552 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 8110 11540 8116 11552
rect 7699 11512 8116 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8536 11512 9137 11540
rect 8536 11500 8542 11512
rect 9125 11509 9137 11512
rect 9171 11540 9183 11543
rect 10888 11540 10916 11580
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 19337 11611 19395 11617
rect 19337 11577 19349 11611
rect 19383 11608 19395 11611
rect 19794 11608 19800 11620
rect 19383 11580 19800 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 19794 11568 19800 11580
rect 19852 11608 19858 11620
rect 20530 11608 20536 11620
rect 19852 11580 20536 11608
rect 19852 11568 19858 11580
rect 20530 11568 20536 11580
rect 20588 11568 20594 11620
rect 16298 11540 16304 11552
rect 9171 11512 10916 11540
rect 16259 11512 16304 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16666 11540 16672 11552
rect 16627 11512 16672 11540
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 20714 11540 20720 11552
rect 20211 11512 20720 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 20714 11500 20720 11512
rect 20772 11540 20778 11552
rect 20990 11540 20996 11552
rect 20772 11512 20996 11540
rect 20772 11500 20778 11512
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2924 11308 3433 11336
rect 2924 11296 2930 11308
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 5626 11336 5632 11348
rect 3467 11308 5632 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9950 11336 9956 11348
rect 9263 11308 9956 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10870 11336 10876 11348
rect 10612 11308 10876 11336
rect 3050 11268 3056 11280
rect 2240 11240 3056 11268
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 2240 11209 2268 11240
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 5353 11271 5411 11277
rect 5353 11237 5365 11271
rect 5399 11268 5411 11271
rect 9398 11268 9404 11280
rect 5399 11240 6132 11268
rect 5399 11237 5411 11240
rect 5353 11231 5411 11237
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 1544 11172 2237 11200
rect 1544 11160 1550 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2225 11163 2283 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 3200 11172 3801 11200
rect 3200 11160 3206 11172
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3789 11163 3847 11169
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5258 11200 5264 11212
rect 4847 11172 5264 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 6104 11209 6132 11240
rect 7300 11240 9404 11268
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6822 11200 6828 11212
rect 6319 11172 6828 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7300 11209 7328 11240
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 10612 11209 10640 11308
rect 10870 11296 10876 11308
rect 10928 11336 10934 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10928 11308 10977 11336
rect 10928 11296 10934 11308
rect 10965 11305 10977 11308
rect 11011 11336 11023 11339
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 11011 11308 11345 11336
rect 11011 11305 11023 11308
rect 10965 11299 11023 11305
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 17218 11336 17224 11348
rect 15519 11308 17224 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 19610 11336 19616 11348
rect 19383 11308 19616 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 10836 11240 13645 11268
rect 10836 11228 10842 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6972 11172 7113 11200
rect 6972 11160 6978 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 10597 11203 10655 11209
rect 8527 11172 9444 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 1394 11092 1400 11144
rect 1452 11132 1458 11144
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1452 11104 2145 11132
rect 1452 11092 1458 11104
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 6932 11132 6960 11160
rect 3568 11104 6960 11132
rect 7009 11135 7067 11141
rect 3568 11092 3574 11104
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 7926 11132 7932 11144
rect 7055 11104 7932 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8662 11132 8668 11144
rect 8343 11104 8668 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 2406 11064 2412 11076
rect 1535 11036 2412 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 4338 11064 4344 11076
rect 4299 11036 4344 11064
rect 4338 11024 4344 11036
rect 4396 11064 4402 11076
rect 4893 11067 4951 11073
rect 4396 11036 4844 11064
rect 4396 11024 4402 11036
rect 1762 10996 1768 11008
rect 1723 10968 1768 10996
rect 1762 10956 1768 10968
rect 1820 10956 1826 11008
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 4816 10996 4844 11036
rect 4893 11033 4905 11067
rect 4939 11064 4951 11067
rect 5442 11064 5448 11076
rect 4939 11036 5448 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5997 11067 6055 11073
rect 5997 11033 6009 11067
rect 6043 11064 6055 11067
rect 7282 11064 7288 11076
rect 6043 11036 7288 11064
rect 6043 11033 6055 11036
rect 5997 11027 6055 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8478 11064 8484 11076
rect 8251 11036 8484 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9416 11064 9444 11172
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 13446 11200 13452 11212
rect 12124 11172 13452 11200
rect 12124 11160 12130 11172
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 13648 11200 13676 11231
rect 13648 11172 14228 11200
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 10330 11135 10388 11141
rect 10330 11132 10342 11135
rect 9548 11104 10342 11132
rect 9548 11092 9554 11104
rect 10330 11101 10342 11104
rect 10376 11101 10388 11135
rect 10330 11095 10388 11101
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13872 11104 14105 11132
rect 13872 11092 13878 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14200 11132 14228 11172
rect 14349 11135 14407 11141
rect 14349 11132 14361 11135
rect 14200 11104 14361 11132
rect 14093 11095 14151 11101
rect 14349 11101 14361 11104
rect 14395 11101 14407 11135
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 14349 11095 14407 11101
rect 15764 11104 16589 11132
rect 9674 11064 9680 11076
rect 9416 11036 9680 11064
rect 9674 11024 9680 11036
rect 9732 11064 9738 11076
rect 10686 11064 10692 11076
rect 9732 11036 10692 11064
rect 9732 11024 9738 11036
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 15764 11008 15792 11104
rect 16577 11101 16589 11104
rect 16623 11132 16635 11135
rect 16666 11132 16672 11144
rect 16623 11104 16672 11132
rect 16623 11101 16635 11104
rect 16577 11095 16635 11101
rect 16666 11092 16672 11104
rect 16724 11132 16730 11144
rect 17862 11132 17868 11144
rect 16724 11104 17868 11132
rect 16724 11092 16730 11104
rect 17862 11092 17868 11104
rect 17920 11132 17926 11144
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17920 11104 18245 11132
rect 17920 11092 17926 11104
rect 18233 11101 18245 11104
rect 18279 11132 18291 11135
rect 18785 11135 18843 11141
rect 18785 11132 18797 11135
rect 18279 11104 18797 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 18785 11101 18797 11104
rect 18831 11101 18843 11135
rect 18785 11095 18843 11101
rect 20622 11092 20628 11144
rect 20680 11132 20686 11144
rect 20717 11135 20775 11141
rect 20717 11132 20729 11135
rect 20680 11104 20729 11132
rect 20680 11092 20686 11104
rect 20717 11101 20729 11104
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 16844 11067 16902 11073
rect 16844 11033 16856 11067
rect 16890 11064 16902 11067
rect 17402 11064 17408 11076
rect 16890 11036 17408 11064
rect 16890 11033 16902 11036
rect 16844 11027 16902 11033
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 19886 11064 19892 11076
rect 17972 11036 19892 11064
rect 4985 10999 5043 11005
rect 4985 10996 4997 10999
rect 2832 10968 2877 10996
rect 4816 10968 4997 10996
rect 2832 10956 2838 10968
rect 4985 10965 4997 10968
rect 5031 10965 5043 10999
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 4985 10959 5043 10965
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6638 10996 6644 11008
rect 6599 10968 6644 10996
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 7834 10996 7840 11008
rect 7795 10968 7840 10996
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 15746 10996 15752 11008
rect 15707 10968 15752 10996
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 17972 11005 18000 11036
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 20472 11067 20530 11073
rect 20472 11033 20484 11067
rect 20518 11064 20530 11067
rect 20806 11064 20812 11076
rect 20518 11036 20812 11064
rect 20518 11033 20530 11036
rect 20472 11027 20530 11033
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 17957 10999 18015 11005
rect 17957 10965 17969 10999
rect 18003 10965 18015 10999
rect 17957 10959 18015 10965
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 2133 10795 2191 10801
rect 2133 10761 2145 10795
rect 2179 10792 2191 10795
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2179 10764 2697 10792
rect 2179 10761 2191 10764
rect 2133 10755 2191 10761
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2924 10764 3065 10792
rect 2924 10752 2930 10764
rect 3053 10761 3065 10764
rect 3099 10792 3111 10795
rect 3418 10792 3424 10804
rect 3099 10764 3424 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 3970 10792 3976 10804
rect 3835 10764 3976 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 2041 10727 2099 10733
rect 2041 10693 2053 10727
rect 2087 10724 2099 10727
rect 2774 10724 2780 10736
rect 2087 10696 2780 10724
rect 2087 10693 2099 10696
rect 2041 10687 2099 10693
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3804 10724 3832 10755
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5994 10792 6000 10804
rect 5031 10764 6000 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6696 10764 6837 10792
rect 6696 10752 6702 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7469 10795 7527 10801
rect 7469 10761 7481 10795
rect 7515 10761 7527 10795
rect 7469 10755 7527 10761
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9306 10792 9312 10804
rect 9263 10764 9312 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 3252 10696 3832 10724
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 3252 10656 3280 10696
rect 5350 10684 5356 10736
rect 5408 10724 5414 10736
rect 7484 10724 7512 10755
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 9416 10764 15056 10792
rect 9416 10724 9444 10764
rect 9950 10724 9956 10736
rect 5408 10696 7512 10724
rect 7576 10696 9444 10724
rect 9508 10696 9956 10724
rect 5408 10684 5414 10696
rect 2464 10628 3280 10656
rect 2464 10616 2470 10628
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 2188 10560 2237 10588
rect 2188 10548 2194 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3252 10597 3280 10628
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5500 10628 5549 10656
rect 5500 10616 5506 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 7576 10656 7604 10696
rect 5537 10619 5595 10625
rect 5644 10628 7604 10656
rect 7837 10659 7895 10665
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 3108 10560 3157 10588
rect 3108 10548 3114 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5644 10588 5672 10628
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 8570 10656 8576 10668
rect 7883 10628 8576 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 6638 10588 6644 10600
rect 5132 10560 5672 10588
rect 6599 10560 6644 10588
rect 5132 10548 5138 10560
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 7282 10588 7288 10600
rect 6779 10560 7288 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7800 10560 7941 10588
rect 7800 10548 7806 10560
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 8159 10560 8493 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8481 10557 8493 10560
rect 8527 10588 8539 10591
rect 9508 10588 9536 10696
rect 9950 10684 9956 10696
rect 10008 10684 10014 10736
rect 12158 10724 12164 10736
rect 10253 10696 12164 10724
rect 10253 10656 10281 10696
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 8527 10560 9536 10588
rect 9600 10628 10281 10656
rect 10341 10659 10399 10665
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 5353 10523 5411 10529
rect 5353 10520 5365 10523
rect 3016 10492 5365 10520
rect 3016 10480 3022 10492
rect 5353 10489 5365 10492
rect 5399 10489 5411 10523
rect 5353 10483 5411 10489
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 8128 10520 8156 10551
rect 6604 10492 8156 10520
rect 6604 10480 6610 10492
rect 8662 10480 8668 10532
rect 8720 10520 8726 10532
rect 9600 10520 9628 10628
rect 10341 10625 10353 10659
rect 10387 10656 10399 10659
rect 10686 10656 10692 10668
rect 10387 10628 10692 10656
rect 10387 10625 10399 10628
rect 10341 10619 10399 10625
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 12434 10656 12440 10668
rect 10744 10628 12440 10656
rect 10744 10616 10750 10628
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 14360 10659 14418 10665
rect 14360 10625 14372 10659
rect 14406 10656 14418 10659
rect 14918 10656 14924 10668
rect 14406 10628 14924 10656
rect 14406 10625 14418 10628
rect 14360 10619 14418 10625
rect 14918 10616 14924 10628
rect 14976 10616 14982 10668
rect 15028 10656 15056 10764
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15252 10764 15485 10792
rect 15252 10752 15258 10764
rect 15473 10761 15485 10764
rect 15519 10792 15531 10795
rect 16022 10792 16028 10804
rect 15519 10764 16028 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17736 10764 19257 10792
rect 17736 10752 17742 10764
rect 19245 10761 19257 10764
rect 19291 10792 19303 10795
rect 19610 10792 19616 10804
rect 19291 10764 19616 10792
rect 19291 10761 19303 10764
rect 19245 10755 19303 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 20680 10764 21189 10792
rect 20680 10752 20686 10764
rect 21177 10761 21189 10764
rect 21223 10761 21235 10795
rect 21177 10755 21235 10761
rect 18046 10684 18052 10736
rect 18104 10733 18110 10736
rect 19794 10733 19800 10736
rect 18104 10727 18168 10733
rect 18104 10693 18122 10727
rect 18156 10693 18168 10727
rect 19788 10724 19800 10733
rect 19755 10696 19800 10724
rect 18104 10687 18168 10693
rect 19788 10687 19800 10696
rect 18104 10684 18110 10687
rect 19794 10684 19800 10687
rect 19852 10684 19858 10736
rect 17126 10656 17132 10668
rect 15028 10628 17132 10656
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 10870 10588 10876 10600
rect 10643 10560 10876 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 10870 10548 10876 10560
rect 10928 10588 10934 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 10928 10560 11529 10588
rect 10928 10548 10934 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 13872 10560 14105 10588
rect 13872 10548 13878 10560
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 19518 10588 19524 10600
rect 19479 10560 19524 10588
rect 14093 10551 14151 10557
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 8720 10492 9628 10520
rect 8720 10480 8726 10492
rect 20806 10480 20812 10532
rect 20864 10520 20870 10532
rect 20901 10523 20959 10529
rect 20901 10520 20913 10523
rect 20864 10492 20913 10520
rect 20864 10480 20870 10492
rect 20901 10489 20913 10492
rect 20947 10489 20959 10523
rect 20901 10483 20959 10489
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4798 10452 4804 10464
rect 4387 10424 4804 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5592 10424 5917 10452
rect 5592 10412 5598 10424
rect 5905 10421 5917 10424
rect 5951 10452 5963 10455
rect 6086 10452 6092 10464
rect 5951 10424 6092 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 7190 10452 7196 10464
rect 7151 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9674 10452 9680 10464
rect 8987 10424 9680 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2866 10248 2872 10260
rect 1627 10220 2872 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 7098 10248 7104 10260
rect 6604 10220 7104 10248
rect 6604 10208 6610 10220
rect 7098 10208 7104 10220
rect 7156 10208 7162 10260
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 9398 10248 9404 10260
rect 8404 10220 9404 10248
rect 2866 10112 2872 10124
rect 2827 10084 2872 10112
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5500 10084 5733 10112
rect 5500 10072 5506 10084
rect 5721 10081 5733 10084
rect 5767 10112 5779 10115
rect 7650 10112 7656 10124
rect 5767 10084 7656 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8404 10112 8432 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10376 10220 10701 10248
rect 10376 10208 10382 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 14458 10248 14464 10260
rect 10689 10211 10747 10217
rect 10796 10220 14464 10248
rect 9968 10180 9996 10208
rect 10796 10180 10824 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 17034 10248 17040 10260
rect 16623 10220 17040 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17954 10248 17960 10260
rect 17144 10220 17960 10248
rect 9968 10152 10824 10180
rect 14550 10140 14556 10192
rect 14608 10180 14614 10192
rect 17144 10180 17172 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 20128 10220 20453 10248
rect 20128 10208 20134 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 20441 10211 20499 10217
rect 14608 10152 17172 10180
rect 14608 10140 14614 10152
rect 16390 10112 16396 10124
rect 7975 10084 8432 10112
rect 11992 10084 16396 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 3418 10044 3424 10056
rect 3331 10016 3424 10044
rect 3418 10004 3424 10016
rect 3476 10044 3482 10056
rect 4706 10044 4712 10056
rect 3476 10016 4712 10044
rect 3476 10004 3482 10016
rect 4706 10004 4712 10016
rect 4764 10044 4770 10056
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4764 10016 4813 10044
rect 4764 10004 4770 10016
rect 4801 10013 4813 10016
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 7742 10044 7748 10056
rect 6687 10016 7748 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10044 9091 10047
rect 9674 10044 9680 10056
rect 9079 10016 9680 10044
rect 9079 10013 9091 10016
rect 9033 10007 9091 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 11992 10044 12020 10084
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 20070 10072 20076 10124
rect 20128 10112 20134 10124
rect 20346 10112 20352 10124
rect 20128 10084 20352 10112
rect 20128 10072 20134 10084
rect 20346 10072 20352 10084
rect 20404 10112 20410 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 20404 10084 21005 10112
rect 20404 10072 20410 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 20993 10075 21051 10081
rect 9784 10016 12020 10044
rect 12069 10047 12127 10053
rect 2041 9979 2099 9985
rect 2041 9945 2053 9979
rect 2087 9976 2099 9979
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 2087 9948 2697 9976
rect 2087 9945 2099 9948
rect 2041 9939 2099 9945
rect 2685 9945 2697 9948
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 8018 9976 8024 9988
rect 7055 9948 8024 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 2314 9908 2320 9920
rect 2275 9880 2320 9908
rect 2314 9868 2320 9880
rect 2372 9868 2378 9920
rect 2777 9911 2835 9917
rect 2777 9877 2789 9911
rect 2823 9908 2835 9911
rect 2958 9908 2964 9920
rect 2823 9880 2964 9908
rect 2823 9877 2835 9880
rect 2777 9871 2835 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 4154 9908 4160 9920
rect 4115 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 7760 9917 7788 9948
rect 8018 9936 8024 9948
rect 8076 9976 8082 9988
rect 9306 9985 9312 9988
rect 9300 9976 9312 9985
rect 8076 9948 8800 9976
rect 9267 9948 9312 9976
rect 8076 9936 8082 9948
rect 4893 9911 4951 9917
rect 4893 9908 4905 9911
rect 4856 9880 4905 9908
rect 4856 9868 4862 9880
rect 4893 9877 4905 9880
rect 4939 9908 4951 9911
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 4939 9880 6193 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 6181 9877 6193 9880
rect 6227 9908 6239 9911
rect 7653 9911 7711 9917
rect 7653 9908 7665 9911
rect 6227 9880 7665 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 7653 9877 7665 9880
rect 7699 9877 7711 9911
rect 7653 9871 7711 9877
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9877 7803 9911
rect 7745 9871 7803 9877
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8570 9908 8576 9920
rect 8435 9880 8576 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8772 9908 8800 9948
rect 9300 9939 9312 9948
rect 9306 9936 9312 9939
rect 9364 9936 9370 9988
rect 9784 9908 9812 10016
rect 12069 10013 12081 10047
rect 12115 10044 12127 10047
rect 13814 10044 13820 10056
rect 12115 10016 13820 10044
rect 12115 10013 12127 10016
rect 12069 10007 12127 10013
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 11802 9979 11860 9985
rect 11802 9976 11814 9979
rect 11204 9948 11814 9976
rect 11204 9936 11210 9948
rect 11802 9945 11814 9948
rect 11848 9945 11860 9979
rect 11802 9939 11860 9945
rect 12452 9920 12480 10016
rect 13814 10004 13820 10016
rect 13872 10044 13878 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13872 10016 14105 10044
rect 13872 10004 13878 10016
rect 14093 10013 14105 10016
rect 14139 10044 14151 10047
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14139 10016 15485 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 15473 10013 15485 10016
rect 15519 10044 15531 10047
rect 15746 10044 15752 10056
rect 15519 10016 15752 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 17920 10016 18613 10044
rect 17920 10004 17926 10016
rect 18601 10013 18613 10016
rect 18647 10044 18659 10047
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 18647 10016 19257 10044
rect 18647 10013 18659 10016
rect 18601 10007 18659 10013
rect 19245 10013 19257 10016
rect 19291 10044 19303 10047
rect 19518 10044 19524 10056
rect 19291 10016 19524 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19518 10004 19524 10016
rect 19576 10044 19582 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19576 10016 19625 10044
rect 19576 10004 19582 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 16942 9976 16948 9988
rect 16855 9948 16948 9976
rect 16942 9936 16948 9948
rect 17000 9976 17006 9988
rect 18334 9979 18392 9985
rect 18334 9976 18346 9979
rect 17000 9948 18346 9976
rect 17000 9936 17006 9948
rect 18334 9945 18346 9948
rect 18380 9945 18392 9979
rect 18334 9939 18392 9945
rect 8772 9880 9812 9908
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10778 9908 10784 9920
rect 10459 9880 10784 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 12434 9908 12440 9920
rect 12395 9880 12440 9908
rect 12434 9868 12440 9880
rect 12492 9868 12498 9920
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 17221 9911 17279 9917
rect 17221 9908 17233 9911
rect 17184 9880 17233 9908
rect 17184 9868 17190 9880
rect 17221 9877 17233 9880
rect 17267 9877 17279 9911
rect 20070 9908 20076 9920
rect 20031 9880 20076 9908
rect 17221 9871 17279 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20622 9868 20628 9920
rect 20680 9908 20686 9920
rect 20809 9911 20867 9917
rect 20809 9908 20821 9911
rect 20680 9880 20821 9908
rect 20680 9868 20686 9880
rect 20809 9877 20821 9880
rect 20855 9877 20867 9911
rect 20809 9871 20867 9877
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 20956 9880 21001 9908
rect 20956 9868 20962 9880
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2924 9676 3188 9704
rect 2924 9664 2930 9676
rect 3160 9648 3188 9676
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 4212 9676 5457 9704
rect 4212 9664 4218 9676
rect 5445 9673 5457 9676
rect 5491 9673 5503 9707
rect 11146 9704 11152 9716
rect 11107 9676 11152 9704
rect 5445 9667 5503 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 14001 9707 14059 9713
rect 14001 9673 14013 9707
rect 14047 9704 14059 9707
rect 14458 9704 14464 9716
rect 14047 9676 14464 9704
rect 14047 9673 14059 9676
rect 14001 9667 14059 9673
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21177 9707 21235 9713
rect 21177 9704 21189 9707
rect 20956 9676 21189 9704
rect 20956 9664 20962 9676
rect 21177 9673 21189 9676
rect 21223 9673 21235 9707
rect 21177 9667 21235 9673
rect 1394 9636 1400 9648
rect 1355 9608 1400 9636
rect 1394 9596 1400 9608
rect 1452 9596 1458 9648
rect 3142 9596 3148 9648
rect 3200 9596 3206 9648
rect 5994 9636 6000 9648
rect 4356 9608 6000 9636
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 4356 9568 4384 9608
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 6420 9608 7389 9636
rect 6420 9596 6426 9608
rect 7377 9605 7389 9608
rect 7423 9636 7435 9639
rect 8202 9636 8208 9648
rect 7423 9608 8208 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 9122 9596 9128 9648
rect 9180 9596 9186 9648
rect 9248 9639 9306 9645
rect 9248 9605 9260 9639
rect 9294 9636 9306 9639
rect 9398 9636 9404 9648
rect 9294 9608 9404 9636
rect 9294 9605 9306 9608
rect 9248 9599 9306 9605
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 10042 9645 10048 9648
rect 10036 9636 10048 9645
rect 10003 9608 10048 9636
rect 10036 9599 10048 9608
rect 10042 9596 10048 9599
rect 10100 9596 10106 9648
rect 10410 9596 10416 9648
rect 10468 9636 10474 9648
rect 10870 9636 10876 9648
rect 10468 9608 10876 9636
rect 10468 9596 10474 9608
rect 10870 9596 10876 9608
rect 10928 9636 10934 9648
rect 12590 9639 12648 9645
rect 12590 9636 12602 9639
rect 10928 9608 12602 9636
rect 10928 9596 10934 9608
rect 12590 9605 12602 9608
rect 12636 9605 12648 9639
rect 12590 9599 12648 9605
rect 16936 9639 16994 9645
rect 16936 9605 16948 9639
rect 16982 9636 16994 9639
rect 17034 9636 17040 9648
rect 16982 9608 17040 9636
rect 16982 9605 16994 9608
rect 16936 9599 16994 9605
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 19460 9639 19518 9645
rect 19460 9605 19472 9639
rect 19506 9636 19518 9639
rect 19610 9636 19616 9648
rect 19506 9608 19616 9636
rect 19506 9605 19518 9608
rect 19460 9599 19518 9605
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 20530 9596 20536 9648
rect 20588 9636 20594 9648
rect 20717 9639 20775 9645
rect 20717 9636 20729 9639
rect 20588 9608 20729 9636
rect 20588 9596 20594 9608
rect 20717 9605 20729 9608
rect 20763 9605 20775 9639
rect 20717 9599 20775 9605
rect 3237 9531 3295 9537
rect 4264 9540 4384 9568
rect 4433 9571 4491 9577
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 2924 9472 2973 9500
rect 2924 9460 2930 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 3108 9472 3157 9500
rect 3108 9460 3114 9472
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 1857 9435 1915 9441
rect 1857 9401 1869 9435
rect 1903 9432 1915 9435
rect 3252 9432 3280 9531
rect 4264 9509 4292 9540
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 4433 9531 4491 9537
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 3602 9432 3608 9444
rect 1903 9404 2636 9432
rect 1903 9401 1915 9404
rect 1857 9395 1915 9401
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2608 9373 2636 9404
rect 2976 9404 3280 9432
rect 3563 9404 3608 9432
rect 2976 9376 3004 9404
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4356 9432 4384 9463
rect 3936 9404 4384 9432
rect 3936 9392 3942 9404
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9364 2651 9367
rect 2958 9364 2964 9376
rect 2639 9336 2964 9364
rect 2639 9333 2651 9336
rect 2593 9327 2651 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 4448 9364 4476 9531
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6086 9568 6092 9580
rect 5776 9540 6092 9568
rect 5776 9528 5782 9540
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6546 9568 6552 9580
rect 6328 9540 6552 9568
rect 6328 9528 6334 9540
rect 6546 9528 6552 9540
rect 6604 9568 6610 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 6604 9540 7297 9568
rect 6604 9528 6610 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 9140 9568 9168 9596
rect 7285 9531 7343 9537
rect 7576 9540 9168 9568
rect 5258 9500 5264 9512
rect 5171 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6730 9500 6736 9512
rect 6288 9472 6736 9500
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 4801 9435 4859 9441
rect 4801 9432 4813 9435
rect 4580 9404 4813 9432
rect 4580 9392 4586 9404
rect 4801 9401 4813 9404
rect 4847 9401 4859 9435
rect 5276 9432 5304 9460
rect 6288 9432 6316 9472
rect 6730 9460 6736 9472
rect 6788 9500 6794 9512
rect 7576 9509 7604 9540
rect 12434 9528 12440 9580
rect 12492 9528 12498 9580
rect 15114 9571 15172 9577
rect 15114 9568 15126 9571
rect 13740 9540 15126 9568
rect 7561 9503 7619 9509
rect 7561 9500 7573 9503
rect 6788 9472 7573 9500
rect 6788 9460 6794 9472
rect 7561 9469 7573 9472
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9500 9551 9503
rect 9674 9500 9680 9512
rect 9539 9472 9680 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9646 9460 9680 9472
rect 9732 9500 9738 9512
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9732 9472 9781 9500
rect 9732 9460 9738 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9500 12403 9503
rect 12452 9500 12480 9528
rect 12391 9472 12480 9500
rect 12391 9469 12403 9472
rect 12345 9463 12403 9469
rect 8113 9435 8171 9441
rect 8113 9432 8125 9435
rect 5276 9404 6316 9432
rect 6748 9404 8125 9432
rect 4801 9395 4859 9401
rect 5902 9364 5908 9376
rect 3292 9336 4476 9364
rect 5863 9336 5908 9364
rect 3292 9324 3298 9336
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6086 9324 6092 9376
rect 6144 9364 6150 9376
rect 6362 9364 6368 9376
rect 6144 9336 6368 9364
rect 6144 9324 6150 9336
rect 6362 9324 6368 9336
rect 6420 9364 6426 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6420 9336 6561 9364
rect 6420 9324 6426 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6748 9364 6776 9404
rect 8113 9401 8125 9404
rect 8159 9432 8171 9435
rect 8478 9432 8484 9444
rect 8159 9404 8484 9432
rect 8159 9401 8171 9404
rect 8113 9395 8171 9401
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 6914 9364 6920 9376
rect 6696 9336 6776 9364
rect 6875 9336 6920 9364
rect 6696 9324 6702 9336
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 9646 9364 9674 9460
rect 11606 9432 11612 9444
rect 11567 9404 11612 9432
rect 11606 9392 11612 9404
rect 11664 9432 11670 9444
rect 12360 9432 12388 9463
rect 11664 9404 12388 9432
rect 11664 9392 11670 9404
rect 9950 9364 9956 9376
rect 9646 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 13740 9373 13768 9540
rect 15114 9537 15126 9540
rect 15160 9537 15172 9571
rect 15114 9531 15172 9537
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15657 9571 15715 9577
rect 15657 9568 15669 9571
rect 15620 9540 15669 9568
rect 15620 9528 15626 9540
rect 15657 9537 15669 9540
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 17954 9568 17960 9580
rect 16448 9540 17960 9568
rect 16448 9528 16454 9540
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 20346 9568 20352 9580
rect 18064 9540 20352 9568
rect 15378 9500 15384 9512
rect 15339 9472 15384 9500
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 15396 9432 15424 9460
rect 16684 9432 16712 9463
rect 18064 9441 18092 9540
rect 20346 9528 20352 9540
rect 20404 9568 20410 9580
rect 20809 9571 20867 9577
rect 20404 9540 20576 9568
rect 20404 9528 20410 9540
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 20548 9509 20576 9540
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 21266 9568 21272 9580
rect 20855 9540 21272 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 19760 9472 19993 9500
rect 19760 9460 19766 9472
rect 19981 9469 19993 9472
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 20533 9503 20591 9509
rect 20533 9469 20545 9503
rect 20579 9469 20591 9503
rect 20533 9463 20591 9469
rect 15396 9404 16712 9432
rect 18049 9435 18107 9441
rect 18049 9401 18061 9435
rect 18095 9401 18107 9435
rect 18049 9395 18107 9401
rect 13725 9367 13783 9373
rect 13725 9364 13737 9367
rect 10560 9336 13737 9364
rect 10560 9324 10566 9336
rect 13725 9333 13737 9336
rect 13771 9333 13783 9367
rect 13725 9327 13783 9333
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 16264 9336 18337 9364
rect 16264 9324 16270 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18325 9327 18383 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1854 9160 1860 9172
rect 1535 9132 1860 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 3292 9132 3341 9160
rect 3292 9120 3298 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5994 9160 6000 9172
rect 4120 9132 6000 9160
rect 4120 9120 4126 9132
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 9766 9160 9772 9172
rect 7340 9132 9772 9160
rect 7340 9120 7346 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10781 9163 10839 9169
rect 10781 9160 10793 9163
rect 10100 9132 10793 9160
rect 10100 9120 10106 9132
rect 10781 9129 10793 9132
rect 10827 9129 10839 9163
rect 10781 9123 10839 9129
rect 12176 9132 13216 9160
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 9306 9092 9312 9104
rect 1452 9064 2774 9092
rect 1452 9052 1458 9064
rect 2746 9024 2774 9064
rect 5460 9064 9312 9092
rect 3326 9024 3332 9036
rect 2746 8996 3332 9024
rect 3326 8984 3332 8996
rect 3384 9024 3390 9036
rect 3878 9024 3884 9036
rect 3384 8996 3884 9024
rect 3384 8984 3390 8996
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 5460 9033 5488 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 5445 9027 5503 9033
rect 4387 8996 5396 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 3050 8956 3056 8968
rect 2823 8928 3056 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4488 8928 4629 8956
rect 4488 8916 4494 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 5368 8956 5396 8996
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5626 9024 5632 9036
rect 5583 8996 5632 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 6880 8996 6925 9024
rect 6880 8984 6886 8996
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 8076 8996 8125 9024
rect 8076 8984 8082 8996
rect 8113 8993 8125 8996
rect 8159 9024 8171 9027
rect 9030 9024 9036 9036
rect 8159 8996 9036 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 11790 9024 11796 9036
rect 10468 8996 11796 9024
rect 10468 8984 10474 8996
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 12176 9024 12204 9132
rect 13188 9092 13216 9132
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13320 9132 13553 9160
rect 13320 9120 13326 9132
rect 13541 9129 13553 9132
rect 13587 9160 13599 9163
rect 13722 9160 13728 9172
rect 13587 9132 13728 9160
rect 13587 9129 13599 9132
rect 13541 9123 13599 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14274 9160 14280 9172
rect 14139 9132 14280 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 17678 9160 17684 9172
rect 14384 9132 17684 9160
rect 14384 9092 14412 9132
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 19610 9120 19616 9172
rect 19668 9160 19674 9172
rect 19668 9132 20944 9160
rect 19668 9120 19674 9132
rect 13188 9064 14412 9092
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 19794 9092 19800 9104
rect 17920 9064 19800 9092
rect 17920 9052 17926 9064
rect 19794 9052 19800 9064
rect 19852 9092 19858 9104
rect 20162 9092 20168 9104
rect 19852 9064 20168 9092
rect 19852 9052 19858 9064
rect 20162 9052 20168 9064
rect 20220 9092 20226 9104
rect 20530 9092 20536 9104
rect 20220 9064 20536 9092
rect 20220 9052 20226 9064
rect 20530 9052 20536 9064
rect 20588 9092 20594 9104
rect 20588 9064 20852 9092
rect 20588 9052 20594 9064
rect 12176 8996 12296 9024
rect 5718 8956 5724 8968
rect 5368 8928 5724 8956
rect 4617 8919 4675 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 5960 8928 6653 8956
rect 5960 8916 5966 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8662 8956 8668 8968
rect 7975 8928 8668 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9950 8956 9956 8968
rect 9447 8928 9956 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9950 8916 9956 8928
rect 10008 8956 10014 8968
rect 10226 8956 10232 8968
rect 10008 8928 10232 8956
rect 10008 8916 10014 8928
rect 10226 8916 10232 8928
rect 10284 8956 10290 8968
rect 10962 8956 10968 8968
rect 10284 8928 10968 8956
rect 10284 8916 10290 8928
rect 10962 8916 10968 8928
rect 11020 8956 11026 8968
rect 11057 8959 11115 8965
rect 11057 8956 11069 8959
rect 11020 8928 11069 8956
rect 11020 8916 11026 8928
rect 11057 8925 11069 8928
rect 11103 8956 11115 8959
rect 11606 8956 11612 8968
rect 11103 8928 11612 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11606 8916 11612 8928
rect 11664 8956 11670 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11664 8928 12173 8956
rect 11664 8916 11670 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 2958 8888 2964 8900
rect 2455 8860 2964 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 6733 8891 6791 8897
rect 5675 8860 6316 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 3234 8820 3240 8832
rect 1452 8792 3240 8820
rect 1452 8780 1458 8792
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5718 8820 5724 8832
rect 5031 8792 5724 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6288 8829 6316 8860
rect 6733 8857 6745 8891
rect 6779 8888 6791 8891
rect 6914 8888 6920 8900
rect 6779 8860 6920 8888
rect 6779 8857 6791 8860
rect 6733 8851 6791 8857
rect 6914 8848 6920 8860
rect 6972 8848 6978 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9646 8891 9704 8897
rect 9646 8888 9658 8891
rect 8536 8860 9658 8888
rect 8536 8848 8542 8860
rect 9646 8857 9658 8860
rect 9692 8857 9704 8891
rect 9646 8851 9704 8857
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 10410 8888 10416 8900
rect 9824 8860 10416 8888
rect 9824 8848 9830 8860
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 12268 8888 12296 8996
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 18782 9024 18788 9036
rect 17092 8996 18788 9024
rect 17092 8984 17098 8996
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 19886 9024 19892 9036
rect 19847 8996 19892 9024
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20824 9033 20852 9064
rect 20916 9033 20944 9132
rect 20809 9027 20867 9033
rect 20809 8993 20821 9027
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 12417 8959 12475 8965
rect 12417 8956 12429 8959
rect 11164 8860 12296 8888
rect 12406 8925 12429 8956
rect 12463 8925 12475 8959
rect 12406 8919 12475 8925
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8789 6331 8823
rect 6273 8783 6331 8789
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6638 8820 6644 8832
rect 6512 8792 6644 8820
rect 6512 8780 6518 8792
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7156 8792 7573 8820
rect 7156 8780 7162 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7708 8792 8033 8820
rect 7708 8780 7714 8792
rect 8021 8789 8033 8792
rect 8067 8820 8079 8823
rect 9033 8823 9091 8829
rect 9033 8820 9045 8823
rect 8067 8792 9045 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 9033 8789 9045 8792
rect 9079 8820 9091 8823
rect 11164 8820 11192 8860
rect 9079 8792 11192 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12406 8820 12434 8919
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 15206 8959 15264 8965
rect 15206 8956 15218 8959
rect 13780 8928 15218 8956
rect 13780 8916 13786 8928
rect 15206 8925 15218 8928
rect 15252 8925 15264 8959
rect 15206 8919 15264 8925
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15436 8928 15485 8956
rect 15436 8916 15442 8928
rect 15473 8925 15485 8928
rect 15519 8956 15531 8959
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15519 8928 15761 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 15749 8925 15761 8928
rect 15795 8956 15807 8959
rect 15838 8956 15844 8968
rect 15795 8928 15844 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16022 8965 16028 8968
rect 16016 8956 16028 8965
rect 15983 8928 16028 8956
rect 16016 8919 16028 8928
rect 16022 8916 16028 8919
rect 16080 8916 16086 8968
rect 19610 8956 19616 8968
rect 18616 8928 19616 8956
rect 13262 8848 13268 8900
rect 13320 8888 13326 8900
rect 15654 8888 15660 8900
rect 13320 8860 15660 8888
rect 13320 8848 13326 8860
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 15856 8888 15884 8916
rect 17497 8891 17555 8897
rect 17497 8888 17509 8891
rect 15856 8860 17509 8888
rect 17497 8857 17509 8860
rect 17543 8888 17555 8891
rect 17954 8888 17960 8900
rect 17543 8860 17960 8888
rect 17543 8857 17555 8860
rect 17497 8851 17555 8857
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 18141 8891 18199 8897
rect 18141 8888 18153 8891
rect 18012 8860 18153 8888
rect 18012 8848 18018 8860
rect 18141 8857 18153 8860
rect 18187 8857 18199 8891
rect 18141 8851 18199 8857
rect 11848 8792 12434 8820
rect 11848 8780 11854 8792
rect 14918 8780 14924 8832
rect 14976 8820 14982 8832
rect 17034 8820 17040 8832
rect 14976 8792 17040 8820
rect 14976 8780 14982 8792
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8820 17187 8823
rect 17218 8820 17224 8832
rect 17175 8792 17224 8820
rect 17175 8789 17187 8792
rect 17129 8783 17187 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17460 8792 17785 8820
rect 17460 8780 17466 8792
rect 17773 8789 17785 8792
rect 17819 8820 17831 8823
rect 18616 8820 18644 8928
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 20254 8956 20260 8968
rect 19843 8928 20260 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 18782 8848 18788 8900
rect 18840 8888 18846 8900
rect 19705 8891 19763 8897
rect 19705 8888 19717 8891
rect 18840 8860 19717 8888
rect 18840 8848 18846 8860
rect 19705 8857 19717 8860
rect 19751 8857 19763 8891
rect 19705 8851 19763 8857
rect 17819 8792 18644 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 18932 8792 19349 8820
rect 18932 8780 18938 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 19337 8783 19395 8789
rect 20349 8823 20407 8829
rect 20349 8789 20361 8823
rect 20395 8820 20407 8823
rect 20530 8820 20536 8832
rect 20395 8792 20536 8820
rect 20395 8789 20407 8792
rect 20349 8783 20407 8789
rect 20530 8780 20536 8792
rect 20588 8780 20594 8832
rect 20717 8823 20775 8829
rect 20717 8789 20729 8823
rect 20763 8820 20775 8823
rect 20806 8820 20812 8832
rect 20763 8792 20812 8820
rect 20763 8789 20775 8792
rect 20717 8783 20775 8789
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1857 8619 1915 8625
rect 1857 8616 1869 8619
rect 1820 8588 1869 8616
rect 1820 8576 1826 8588
rect 1857 8585 1869 8588
rect 1903 8585 1915 8619
rect 1857 8579 1915 8585
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2004 8588 2329 8616
rect 2004 8576 2010 8588
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 4522 8616 4528 8628
rect 4483 8588 4528 8616
rect 2317 8579 2375 8585
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5534 8616 5540 8628
rect 4948 8588 5028 8616
rect 5495 8588 5540 8616
rect 4948 8576 4954 8588
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 5000 8557 5028 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7892 8588 8033 8616
rect 7892 8576 7898 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8202 8616 8208 8628
rect 8159 8588 8208 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 15102 8616 15108 8628
rect 8312 8588 15108 8616
rect 4985 8551 5043 8557
rect 2924 8520 3832 8548
rect 2924 8508 2930 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8381 1823 8415
rect 1765 8375 1823 8381
rect 2777 8415 2835 8421
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 2866 8412 2872 8424
rect 2823 8384 2872 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 1780 8344 1808 8375
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 3804 8421 3832 8520
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 5031 8520 7021 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 7009 8517 7021 8520
rect 7055 8548 7067 8551
rect 8312 8548 8340 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 16761 8619 16819 8625
rect 16761 8616 16773 8619
rect 15304 8588 16773 8616
rect 7055 8520 8340 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 8720 8520 9137 8548
rect 8720 8508 8726 8520
rect 9125 8517 9137 8520
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 14918 8548 14924 8560
rect 9548 8520 14924 8548
rect 9548 8508 9554 8520
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 4246 8480 4252 8492
rect 4159 8452 4252 8480
rect 4246 8440 4252 8452
rect 4304 8480 4310 8492
rect 4706 8480 4712 8492
rect 4304 8452 4712 8480
rect 4304 8440 4310 8452
rect 4706 8440 4712 8452
rect 4764 8480 4770 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4764 8452 4905 8480
rect 4764 8440 4770 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 6914 8480 6920 8492
rect 4893 8443 4951 8449
rect 5000 8452 6920 8480
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 5000 8412 5028 8452
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 14458 8480 14464 8492
rect 8536 8452 14464 8480
rect 8536 8440 8542 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 15217 8483 15275 8489
rect 15217 8449 15229 8483
rect 15263 8480 15275 8483
rect 15304 8480 15332 8588
rect 16761 8585 16773 8588
rect 16807 8616 16819 8619
rect 17126 8616 17132 8628
rect 16807 8588 17132 8616
rect 16807 8585 16819 8588
rect 16761 8579 16819 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18966 8576 18972 8628
rect 19024 8616 19030 8628
rect 19024 8588 19472 8616
rect 19024 8576 19030 8588
rect 19058 8508 19064 8560
rect 19116 8548 19122 8560
rect 19254 8551 19312 8557
rect 19254 8548 19266 8551
rect 19116 8520 19266 8548
rect 19116 8508 19122 8520
rect 19254 8517 19266 8520
rect 19300 8517 19312 8551
rect 19254 8511 19312 8517
rect 15263 8452 15332 8480
rect 15263 8449 15275 8452
rect 15217 8443 15275 8449
rect 3835 8384 5028 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 5074 8372 5080 8424
rect 5132 8412 5138 8424
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 5132 8384 5181 8412
rect 5132 8372 5138 8384
rect 5169 8381 5181 8384
rect 5215 8412 5227 8415
rect 5258 8412 5264 8424
rect 5215 8384 5264 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 7282 8412 7288 8424
rect 6380 8384 7288 8412
rect 2130 8344 2136 8356
rect 1780 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8344 2194 8356
rect 3237 8347 3295 8353
rect 3237 8344 3249 8347
rect 2188 8316 3249 8344
rect 2188 8304 2194 8316
rect 3237 8313 3249 8316
rect 3283 8344 3295 8347
rect 6380 8344 6408 8384
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 7975 8384 8892 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 6546 8344 6552 8356
rect 3283 8316 6408 8344
rect 6507 8316 6552 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 8478 8276 8484 8288
rect 8439 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8754 8276 8760 8288
rect 8715 8248 8760 8276
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 8864 8276 8892 8384
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 13262 8412 13268 8424
rect 9272 8384 13268 8412
rect 9272 8372 9278 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 14274 8412 14280 8424
rect 13412 8384 14280 8412
rect 13412 8372 13418 8384
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15838 8412 15844 8424
rect 15519 8384 15844 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 19444 8412 19472 8588
rect 19720 8520 21220 8548
rect 19720 8492 19748 8520
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19702 8480 19708 8492
rect 19567 8452 19708 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 21192 8489 21220 8520
rect 20910 8483 20968 8489
rect 20910 8480 20922 8483
rect 19996 8452 20922 8480
rect 19996 8412 20024 8452
rect 20910 8449 20922 8452
rect 20956 8449 20968 8483
rect 20910 8443 20968 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 19444 8384 20024 8412
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 11790 8344 11796 8356
rect 9088 8316 11796 8344
rect 9088 8304 9094 8316
rect 11790 8304 11796 8316
rect 11848 8344 11854 8356
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 11848 8316 14105 8344
rect 11848 8304 11854 8316
rect 14093 8313 14105 8316
rect 14139 8313 14151 8347
rect 18230 8344 18236 8356
rect 14093 8307 14151 8313
rect 15488 8316 18236 8344
rect 9214 8276 9220 8288
rect 8864 8248 9220 8276
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9677 8279 9735 8285
rect 9677 8245 9689 8279
rect 9723 8276 9735 8279
rect 10226 8276 10232 8288
rect 9723 8248 10232 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 10226 8236 10232 8248
rect 10284 8276 10290 8288
rect 10413 8279 10471 8285
rect 10413 8276 10425 8279
rect 10284 8248 10425 8276
rect 10284 8236 10290 8248
rect 10413 8245 10425 8248
rect 10459 8245 10471 8279
rect 10413 8239 10471 8245
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 12158 8276 12164 8288
rect 10652 8248 12164 8276
rect 10652 8236 10658 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 13630 8276 13636 8288
rect 13591 8248 13636 8276
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15488 8276 15516 8316
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19794 8344 19800 8356
rect 19755 8316 19800 8344
rect 19794 8304 19800 8316
rect 19852 8304 19858 8356
rect 15838 8276 15844 8288
rect 15160 8248 15516 8276
rect 15799 8248 15844 8276
rect 15160 8236 15166 8248
rect 15838 8236 15844 8248
rect 15896 8276 15902 8288
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 15896 8248 16129 8276
rect 15896 8236 15902 8248
rect 16117 8245 16129 8248
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 16390 8236 16396 8288
rect 16448 8276 16454 8288
rect 17402 8276 17408 8288
rect 16448 8248 17408 8276
rect 16448 8236 16454 8248
rect 17402 8236 17408 8248
rect 17460 8276 17466 8288
rect 18141 8279 18199 8285
rect 18141 8276 18153 8279
rect 17460 8248 18153 8276
rect 17460 8236 17466 8248
rect 18141 8245 18153 8248
rect 18187 8245 18199 8279
rect 18141 8239 18199 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 3970 8072 3976 8084
rect 2464 8044 3976 8072
rect 2464 8032 2470 8044
rect 3970 8032 3976 8044
rect 4028 8072 4034 8084
rect 4157 8075 4215 8081
rect 4157 8072 4169 8075
rect 4028 8044 4169 8072
rect 4028 8032 4034 8044
rect 4157 8041 4169 8044
rect 4203 8041 4215 8075
rect 4157 8035 4215 8041
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5994 8072 6000 8084
rect 5132 8044 6000 8072
rect 5132 8032 5138 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9582 8072 9588 8084
rect 8987 8044 9588 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 12158 8032 12164 8084
rect 12216 8072 12222 8084
rect 17954 8072 17960 8084
rect 12216 8044 17172 8072
rect 17915 8044 17960 8072
rect 12216 8032 12222 8044
rect 3142 8004 3148 8016
rect 1780 7976 3148 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1780 7945 1808 7976
rect 3142 7964 3148 7976
rect 3200 8004 3206 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3200 7976 3801 8004
rect 3200 7964 3206 7976
rect 3789 7973 3801 7976
rect 3835 8004 3847 8007
rect 4062 8004 4068 8016
rect 3835 7976 4068 8004
rect 3835 7973 3847 7976
rect 3789 7967 3847 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 6546 8004 6552 8016
rect 5460 7976 6552 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7905 1823 7939
rect 1765 7899 1823 7905
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7936 2743 7939
rect 2731 7908 3188 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 1688 7868 1716 7896
rect 2406 7868 2412 7880
rect 1688 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 1578 7760 1584 7812
rect 1636 7800 1642 7812
rect 2777 7803 2835 7809
rect 2777 7800 2789 7803
rect 1636 7772 2789 7800
rect 1636 7760 1642 7772
rect 2777 7769 2789 7772
rect 2823 7769 2835 7803
rect 3160 7800 3188 7908
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 5460 7936 5488 7976
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 7064 7976 8248 8004
rect 7064 7964 7070 7976
rect 8220 7948 8248 7976
rect 4028 7908 5488 7936
rect 5537 7939 5595 7945
rect 4028 7896 4034 7908
rect 5537 7905 5549 7939
rect 5583 7905 5595 7939
rect 5718 7936 5724 7948
rect 5679 7908 5724 7936
rect 5537 7899 5595 7905
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 3510 7868 3516 7880
rect 3292 7840 3516 7868
rect 3292 7828 3298 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 5552 7868 5580 7899
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7098 7936 7104 7948
rect 7059 7908 7104 7936
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 15838 7936 15844 7948
rect 15344 7908 15844 7936
rect 15344 7896 15350 7908
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 17144 7936 17172 8044
rect 17954 8032 17960 8044
rect 18012 8072 18018 8084
rect 18322 8072 18328 8084
rect 18012 8044 18328 8072
rect 18012 8032 18018 8044
rect 18322 8032 18328 8044
rect 18380 8072 18386 8084
rect 18785 8075 18843 8081
rect 18785 8072 18797 8075
rect 18380 8044 18797 8072
rect 18380 8032 18386 8044
rect 18785 8041 18797 8044
rect 18831 8041 18843 8075
rect 18785 8035 18843 8041
rect 19981 8075 20039 8081
rect 19981 8041 19993 8075
rect 20027 8072 20039 8075
rect 20438 8072 20444 8084
rect 20027 8044 20444 8072
rect 20027 8041 20039 8044
rect 19981 8035 20039 8041
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 20990 8072 20996 8084
rect 20951 8044 20996 8072
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 17221 8007 17279 8013
rect 17221 7973 17233 8007
rect 17267 8004 17279 8007
rect 19058 8004 19064 8016
rect 17267 7976 19064 8004
rect 17267 7973 17279 7976
rect 17221 7967 17279 7973
rect 19058 7964 19064 7976
rect 19116 8004 19122 8016
rect 19116 7976 19380 8004
rect 19116 7964 19122 7976
rect 18046 7936 18052 7948
rect 17144 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 19352 7945 19380 7976
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 21269 8007 21327 8013
rect 21269 8004 21281 8007
rect 20312 7976 21281 8004
rect 20312 7964 20318 7976
rect 21269 7973 21281 7976
rect 21315 7973 21327 8007
rect 21269 7967 21327 7973
rect 19337 7939 19395 7945
rect 19337 7905 19349 7939
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7905 20407 7939
rect 20530 7936 20536 7948
rect 20491 7908 20536 7936
rect 20349 7899 20407 7905
rect 9214 7868 9220 7880
rect 5552 7840 9220 7868
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 10054 7871 10112 7877
rect 10054 7868 10066 7871
rect 9364 7840 10066 7868
rect 9364 7828 9370 7840
rect 10054 7837 10066 7840
rect 10100 7868 10112 7871
rect 10100 7840 10180 7868
rect 10100 7837 10112 7840
rect 10054 7831 10112 7837
rect 3160 7772 3372 7800
rect 2777 7763 2835 7769
rect 1854 7732 1860 7744
rect 1815 7704 1860 7732
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3344 7732 3372 7772
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 8021 7803 8079 7809
rect 3476 7772 6684 7800
rect 3476 7760 3482 7772
rect 5258 7732 5264 7744
rect 3344 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7732 5322 7744
rect 5718 7732 5724 7744
rect 5316 7704 5724 7732
rect 5316 7692 5322 7704
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5994 7732 6000 7744
rect 5859 7704 6000 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6546 7732 6552 7744
rect 6227 7704 6552 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6656 7741 6684 7772
rect 8021 7769 8033 7803
rect 8067 7800 8079 7803
rect 8662 7800 8668 7812
rect 8067 7772 8668 7800
rect 8067 7769 8079 7772
rect 8021 7763 8079 7769
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 6641 7735 6699 7741
rect 6641 7701 6653 7735
rect 6687 7701 6699 7735
rect 7006 7732 7012 7744
rect 6967 7704 7012 7732
rect 6641 7695 6699 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8478 7732 8484 7744
rect 8159 7704 8484 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 10152 7732 10180 7840
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10284 7840 10333 7868
rect 10284 7828 10290 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10336 7800 10364 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11710 7871 11768 7877
rect 11710 7868 11722 7871
rect 11204 7840 11722 7868
rect 11204 7828 11210 7840
rect 11710 7837 11722 7840
rect 11756 7837 11768 7871
rect 11710 7831 11768 7837
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 10336 7772 11744 7800
rect 11716 7744 11744 7772
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10152 7704 10609 7732
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 11992 7732 12020 7831
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 16114 7877 16120 7880
rect 16097 7871 16120 7877
rect 16097 7868 16109 7871
rect 15712 7840 16109 7868
rect 15712 7828 15718 7840
rect 16097 7837 16109 7840
rect 16172 7868 16178 7880
rect 16172 7840 16245 7868
rect 16097 7831 16120 7837
rect 16114 7828 16120 7831
rect 16172 7828 16178 7840
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 17460 7840 19533 7868
rect 17460 7828 17466 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 20254 7868 20260 7880
rect 20036 7840 20260 7868
rect 20036 7828 20042 7840
rect 20254 7828 20260 7840
rect 20312 7868 20318 7880
rect 20364 7868 20392 7899
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 20312 7840 20392 7868
rect 20312 7828 20318 7840
rect 14458 7760 14464 7812
rect 14516 7800 14522 7812
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 14516 7772 19625 7800
rect 14516 7760 14522 7772
rect 19613 7769 19625 7772
rect 19659 7769 19671 7803
rect 19613 7763 19671 7769
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 11756 7704 12265 7732
rect 11756 7692 11762 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 17310 7692 17316 7744
rect 17368 7732 17374 7744
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17368 7704 17509 7732
rect 17368 7692 17374 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 19978 7732 19984 7744
rect 18555 7704 19984 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20438 7692 20444 7744
rect 20496 7732 20502 7744
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 20496 7704 20637 7732
rect 20496 7692 20502 7704
rect 20625 7701 20637 7704
rect 20671 7701 20683 7735
rect 20625 7695 20683 7701
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3375 7500 3985 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4120 7500 4353 7528
rect 4120 7488 4126 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4890 7528 4896 7540
rect 4479 7500 4896 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 5994 7528 6000 7540
rect 5955 7500 6000 7528
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8260 7500 8953 7528
rect 8260 7488 8266 7500
rect 8941 7497 8953 7500
rect 8987 7528 8999 7531
rect 10778 7528 10784 7540
rect 8987 7500 10784 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 17586 7528 17592 7540
rect 16715 7500 17592 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 19475 7500 20177 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 20165 7497 20177 7500
rect 20211 7497 20223 7531
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 20165 7491 20223 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 5629 7463 5687 7469
rect 5629 7460 5641 7463
rect 3292 7432 5641 7460
rect 3292 7420 3298 7432
rect 5629 7429 5641 7432
rect 5675 7429 5687 7463
rect 7282 7460 7288 7472
rect 5629 7423 5687 7429
rect 5736 7432 7288 7460
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 5736 7392 5764 7432
rect 7282 7420 7288 7432
rect 7340 7460 7346 7472
rect 10594 7460 10600 7472
rect 7340 7432 10600 7460
rect 7340 7420 7346 7432
rect 10594 7420 10600 7432
rect 10652 7420 10658 7472
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 10744 7432 13943 7460
rect 10744 7420 10750 7432
rect 4632 7364 5764 7392
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2041 7287 2099 7293
rect 2056 7256 2084 7287
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2774 7324 2780 7336
rect 2740 7296 2780 7324
rect 2740 7284 2746 7296
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 3970 7324 3976 7336
rect 3651 7296 3976 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 3620 7256 3648 7287
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4632 7333 4660 7364
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7248 7364 7941 7392
rect 7248 7352 7254 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 10514 7395 10572 7401
rect 10514 7392 10526 7395
rect 9272 7364 10526 7392
rect 9272 7352 9278 7364
rect 10514 7361 10526 7364
rect 10560 7361 10572 7395
rect 10514 7355 10572 7361
rect 12641 7395 12699 7401
rect 12641 7361 12653 7395
rect 12687 7392 12699 7395
rect 13446 7392 13452 7404
rect 12687 7364 13452 7392
rect 12687 7361 12699 7364
rect 12641 7355 12699 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13915 7401 13943 7432
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 21284 7460 21312 7488
rect 19024 7432 21312 7460
rect 19024 7420 19030 7432
rect 13900 7395 13958 7401
rect 13900 7361 13912 7395
rect 13946 7392 13958 7395
rect 17793 7395 17851 7401
rect 13946 7364 15792 7392
rect 13946 7361 13958 7364
rect 13900 7355 13958 7361
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 4120 7296 4629 7324
rect 4120 7284 4126 7296
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5353 7287 5411 7293
rect 2056 7228 3648 7256
rect 5368 7256 5396 7287
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 8202 7324 8208 7336
rect 8163 7296 8208 7324
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 12943 7296 13645 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 5626 7256 5632 7268
rect 5368 7228 5632 7256
rect 5626 7216 5632 7228
rect 5684 7256 5690 7268
rect 9766 7256 9772 7268
rect 5684 7228 9772 7256
rect 5684 7216 5690 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7558 7188 7564 7200
rect 7331 7160 7564 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 7653 7191 7711 7197
rect 7653 7157 7665 7191
rect 7699 7188 7711 7191
rect 7834 7188 7840 7200
rect 7699 7160 7840 7188
rect 7699 7157 7711 7160
rect 7653 7151 7711 7157
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 9180 7160 9413 7188
rect 9180 7148 9186 7160
rect 9401 7157 9413 7160
rect 9447 7188 9459 7191
rect 10042 7188 10048 7200
rect 9447 7160 10048 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10796 7188 10824 7287
rect 11054 7188 11060 7200
rect 10796 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 13280 7197 13308 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 15286 7256 15292 7268
rect 14568 7228 15292 7256
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11204 7160 11529 7188
rect 11204 7148 11210 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13630 7188 13636 7200
rect 13311 7160 13636 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13630 7148 13636 7160
rect 13688 7188 13694 7200
rect 14568 7188 14596 7228
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 15764 7265 15792 7364
rect 17793 7361 17805 7395
rect 17839 7392 17851 7395
rect 17954 7392 17960 7404
rect 17839 7364 17960 7392
rect 17839 7361 17851 7364
rect 17793 7355 17851 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7392 18107 7395
rect 18322 7392 18328 7404
rect 18095 7364 18328 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 20530 7392 20536 7404
rect 20491 7364 20536 7392
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7392 20683 7395
rect 21174 7392 21180 7404
rect 20671 7364 21180 7392
rect 20671 7361 20683 7364
rect 20625 7355 20683 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 17972 7324 18000 7352
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 17972 7296 18705 7324
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19337 7327 19395 7333
rect 19337 7324 19349 7327
rect 19116 7296 19349 7324
rect 19116 7284 19122 7296
rect 19337 7293 19349 7296
rect 19383 7324 19395 7327
rect 20070 7324 20076 7336
rect 19383 7296 20076 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 20717 7327 20775 7333
rect 20717 7293 20729 7327
rect 20763 7293 20775 7327
rect 20717 7287 20775 7293
rect 15749 7259 15807 7265
rect 15749 7225 15761 7259
rect 15795 7256 15807 7259
rect 16298 7256 16304 7268
rect 15795 7228 16304 7256
rect 15795 7225 15807 7228
rect 15749 7219 15807 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 18414 7216 18420 7268
rect 18472 7256 18478 7268
rect 19889 7259 19947 7265
rect 19889 7256 19901 7259
rect 18472 7228 19901 7256
rect 18472 7216 18478 7228
rect 19889 7225 19901 7228
rect 19935 7225 19947 7259
rect 19889 7219 19947 7225
rect 20346 7216 20352 7268
rect 20404 7256 20410 7268
rect 20732 7256 20760 7287
rect 20404 7228 20760 7256
rect 20404 7216 20410 7228
rect 15010 7188 15016 7200
rect 13688 7160 14596 7188
rect 14971 7160 15016 7188
rect 13688 7148 13694 7160
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 15620 7160 16221 7188
rect 15620 7148 15626 7160
rect 16209 7157 16221 7160
rect 16255 7188 16267 7191
rect 16390 7188 16396 7200
rect 16255 7160 16396 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2280 6956 2421 6984
rect 2280 6944 2286 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7064 6956 7481 6984
rect 7064 6944 7070 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 7469 6947 7527 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9324 6956 15792 6984
rect 3418 6916 3424 6928
rect 3068 6888 3424 6916
rect 3068 6857 3096 6888
rect 3418 6876 3424 6888
rect 3476 6916 3482 6928
rect 4062 6916 4068 6928
rect 3476 6888 4068 6916
rect 3476 6876 3482 6888
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 7558 6916 7564 6928
rect 4816 6888 5856 6916
rect 4816 6857 4844 6888
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6817 3111 6851
rect 3053 6811 3111 6817
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5828 6857 5856 6888
rect 6656 6888 7564 6916
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5132 6820 5641 6848
rect 5132 6808 5138 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5994 6848 6000 6860
rect 5859 6820 6000 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6656 6857 6684 6888
rect 7558 6876 7564 6888
rect 7616 6916 7622 6928
rect 9324 6916 9352 6956
rect 7616 6888 9352 6916
rect 12069 6919 12127 6925
rect 7616 6876 7622 6888
rect 12069 6885 12081 6919
rect 12115 6885 12127 6919
rect 15764 6916 15792 6956
rect 18414 6944 18420 6996
rect 18472 6984 18478 6996
rect 19058 6984 19064 6996
rect 18472 6956 19064 6984
rect 18472 6944 18478 6956
rect 19058 6944 19064 6956
rect 19116 6944 19122 6996
rect 17954 6916 17960 6928
rect 15764 6888 17960 6916
rect 12069 6879 12127 6885
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7929 6851 7987 6857
rect 7929 6848 7941 6851
rect 6880 6820 7941 6848
rect 6880 6808 6886 6820
rect 7929 6817 7941 6820
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 12084 6848 12112 6879
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18322 6876 18328 6928
rect 18380 6916 18386 6928
rect 18598 6916 18604 6928
rect 18380 6888 18604 6916
rect 18380 6876 18386 6888
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 8076 6820 8121 6848
rect 10520 6820 12112 6848
rect 17589 6851 17647 6857
rect 8076 6808 8082 6820
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 3142 6780 3148 6792
rect 1535 6752 3148 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 3142 6740 3148 6752
rect 3200 6780 3206 6792
rect 3418 6780 3424 6792
rect 3200 6752 3424 6780
rect 3200 6740 3206 6752
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 4890 6780 4896 6792
rect 4663 6752 4896 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4890 6740 4896 6752
rect 4948 6780 4954 6792
rect 5350 6780 5356 6792
rect 4948 6752 5356 6780
rect 4948 6740 4954 6752
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 6914 6780 6920 6792
rect 6779 6752 6920 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7466 6780 7472 6792
rect 7156 6752 7472 6780
rect 7156 6740 7162 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10330 6783 10388 6789
rect 10330 6780 10342 6783
rect 9824 6752 10342 6780
rect 9824 6740 9830 6752
rect 10330 6749 10342 6752
rect 10376 6780 10388 6783
rect 10520 6780 10548 6820
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 20070 6848 20076 6860
rect 17635 6820 20076 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20404 6820 21189 6848
rect 20404 6808 20410 6820
rect 21177 6817 21189 6820
rect 21223 6817 21235 6851
rect 21177 6811 21235 6817
rect 10376 6752 10548 6780
rect 10597 6783 10655 6789
rect 10376 6749 10388 6752
rect 10330 6743 10388 6749
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 11054 6780 11060 6792
rect 10643 6752 11060 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11974 6780 11980 6792
rect 11164 6752 11980 6780
rect 1762 6672 1768 6724
rect 1820 6712 1826 6724
rect 2777 6715 2835 6721
rect 2777 6712 2789 6715
rect 1820 6684 2789 6712
rect 1820 6672 1826 6684
rect 2777 6681 2789 6684
rect 2823 6681 2835 6715
rect 5537 6715 5595 6721
rect 5537 6712 5549 6715
rect 2777 6675 2835 6681
rect 3804 6684 5549 6712
rect 3804 6656 3832 6684
rect 5537 6681 5549 6684
rect 5583 6681 5595 6715
rect 5537 6675 5595 6681
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 5868 6684 7236 6712
rect 5868 6672 5874 6684
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2179 6616 2881 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2869 6613 2881 6616
rect 2915 6644 2927 6647
rect 3050 6644 3056 6656
rect 2915 6616 3056 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3050 6604 3056 6616
rect 3108 6644 3114 6656
rect 3234 6644 3240 6656
rect 3108 6616 3240 6644
rect 3108 6604 3114 6616
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4522 6644 4528 6656
rect 4483 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 7006 6644 7012 6656
rect 6871 6616 7012 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7208 6653 7236 6684
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 8536 6684 8585 6712
rect 8536 6672 8542 6684
rect 8573 6681 8585 6684
rect 8619 6712 8631 6715
rect 10502 6712 10508 6724
rect 8619 6684 10508 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 10502 6672 10508 6684
rect 10560 6712 10566 6724
rect 11164 6712 11192 6752
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13630 6780 13636 6792
rect 13495 6752 13636 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13688 6752 14105 6780
rect 13688 6740 13694 6752
rect 14093 6749 14105 6752
rect 14139 6780 14151 6783
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14139 6752 14565 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14553 6749 14565 6752
rect 14599 6780 14611 6783
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 14599 6752 16221 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 16209 6749 16221 6752
rect 16255 6749 16267 6783
rect 17310 6780 17316 6792
rect 17271 6752 17316 6780
rect 16209 6743 16267 6749
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6780 17463 6783
rect 18874 6780 18880 6792
rect 17451 6752 18880 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 20162 6780 20168 6792
rect 20027 6752 20168 6780
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 10560 6684 11192 6712
rect 10560 6672 10566 6684
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 13182 6715 13240 6721
rect 13182 6712 13194 6715
rect 11296 6684 13194 6712
rect 11296 6672 11302 6684
rect 13182 6681 13194 6684
rect 13228 6681 13240 6715
rect 13182 6675 13240 6681
rect 14820 6715 14878 6721
rect 14820 6681 14832 6715
rect 14866 6712 14878 6715
rect 16022 6712 16028 6724
rect 14866 6684 16028 6712
rect 14866 6681 14878 6684
rect 14820 6675 14878 6681
rect 16022 6672 16028 6684
rect 16080 6712 16086 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16080 6684 16681 6712
rect 16080 6672 16086 6684
rect 16669 6681 16681 6684
rect 16715 6712 16727 6715
rect 18506 6712 18512 6724
rect 16715 6684 18512 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 18782 6712 18788 6724
rect 18743 6684 18788 6712
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 20349 6715 20407 6721
rect 20349 6681 20361 6715
rect 20395 6712 20407 6715
rect 20806 6712 20812 6724
rect 20395 6684 20812 6712
rect 20395 6681 20407 6684
rect 20349 6675 20407 6681
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6613 7251 6647
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7193 6607 7251 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9398 6644 9404 6656
rect 9180 6616 9404 6644
rect 9180 6604 9186 6616
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11054 6644 11060 6656
rect 11011 6616 11060 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11698 6644 11704 6656
rect 11112 6616 11704 6644
rect 11112 6604 11118 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 15933 6647 15991 6653
rect 15933 6644 15945 6647
rect 15804 6616 15945 6644
rect 15804 6604 15810 6616
rect 15933 6613 15945 6616
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 16945 6647 17003 6653
rect 16945 6613 16957 6647
rect 16991 6644 17003 6647
rect 17126 6644 17132 6656
rect 16991 6616 17132 6644
rect 16991 6613 17003 6616
rect 16945 6607 17003 6613
rect 17126 6604 17132 6616
rect 17184 6604 17190 6656
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6644 18199 6647
rect 18230 6644 18236 6656
rect 18187 6616 18236 6644
rect 18187 6613 18199 6616
rect 18141 6607 18199 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 18414 6644 18420 6656
rect 18375 6616 18420 6644
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 18598 6604 18604 6656
rect 18656 6644 18662 6656
rect 19337 6647 19395 6653
rect 19337 6644 19349 6647
rect 18656 6616 19349 6644
rect 18656 6604 18662 6616
rect 19337 6613 19349 6616
rect 19383 6644 19395 6647
rect 19518 6644 19524 6656
rect 19383 6616 19524 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 19610 6604 19616 6656
rect 19668 6644 19674 6656
rect 20364 6644 20392 6675
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 20993 6715 21051 6721
rect 20993 6681 21005 6715
rect 21039 6712 21051 6715
rect 21358 6712 21364 6724
rect 21039 6684 21364 6712
rect 21039 6681 21051 6684
rect 20993 6675 21051 6681
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 20622 6644 20628 6656
rect 19668 6616 20392 6644
rect 20583 6616 20628 6644
rect 19668 6604 19674 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20898 6604 20904 6656
rect 20956 6644 20962 6656
rect 21085 6647 21143 6653
rect 21085 6644 21097 6647
rect 20956 6616 21097 6644
rect 20956 6604 20962 6616
rect 21085 6613 21097 6616
rect 21131 6613 21143 6647
rect 21085 6607 21143 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1946 6440 1952 6452
rect 1627 6412 1952 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2590 6440 2596 6452
rect 2551 6412 2596 6440
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 3016 6412 3065 6440
rect 3016 6400 3022 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 4890 6440 4896 6452
rect 4851 6412 4896 6440
rect 3053 6403 3111 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5316 6412 5733 6440
rect 5316 6400 5322 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 7929 6443 7987 6449
rect 7929 6409 7941 6443
rect 7975 6440 7987 6443
rect 9582 6440 9588 6452
rect 7975 6412 9588 6440
rect 7975 6409 7987 6412
rect 7929 6403 7987 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 13446 6440 13452 6452
rect 13407 6412 13452 6440
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 16301 6443 16359 6449
rect 16301 6440 16313 6443
rect 15528 6412 16313 6440
rect 15528 6400 15534 6412
rect 16301 6409 16313 6412
rect 16347 6409 16359 6443
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 16301 6403 16359 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18969 6443 19027 6449
rect 18969 6440 18981 6443
rect 18012 6412 18981 6440
rect 18012 6400 18018 6412
rect 18969 6409 18981 6412
rect 19015 6409 19027 6443
rect 18969 6403 19027 6409
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 7064 6344 7604 6372
rect 7064 6332 7070 6344
rect 7576 6316 7604 6344
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 8481 6375 8539 6381
rect 8481 6372 8493 6375
rect 7800 6344 8493 6372
rect 7800 6332 7806 6344
rect 8481 6341 8493 6344
rect 8527 6341 8539 6375
rect 8481 6335 8539 6341
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 15930 6372 15936 6384
rect 8904 6344 12204 6372
rect 15891 6344 15936 6372
rect 8904 6332 8910 6344
rect 12176 6316 12204 6344
rect 15930 6332 15936 6344
rect 15988 6332 15994 6384
rect 18693 6375 18751 6381
rect 16040 6344 18184 6372
rect 1394 6264 1400 6316
rect 1452 6304 1458 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1452 6276 1961 6304
rect 1452 6264 1458 6276
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2740 6276 2973 6304
rect 2740 6264 2746 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 4246 6304 4252 6316
rect 4159 6276 4252 6304
rect 2961 6267 3019 6273
rect 4246 6264 4252 6276
rect 4304 6304 4310 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 4304 6276 5641 6304
rect 4304 6264 4310 6276
rect 5629 6273 5641 6276
rect 5675 6304 5687 6307
rect 6914 6304 6920 6316
rect 5675 6276 6132 6304
rect 6827 6276 6920 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 1820 6208 2053 6236
rect 1820 6196 1826 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2314 6236 2320 6248
rect 2271 6208 2320 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 1578 6128 1584 6180
rect 1636 6168 1642 6180
rect 2240 6168 2268 6199
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3970 6236 3976 6248
rect 3283 6208 3976 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5905 6239 5963 6245
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 5994 6236 6000 6248
rect 5951 6208 6000 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6104 6236 6132 6276
rect 6914 6264 6920 6276
rect 6972 6304 6978 6316
rect 6972 6276 7512 6304
rect 6972 6264 6978 6276
rect 7484 6248 7512 6276
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8570 6304 8576 6316
rect 7616 6276 7661 6304
rect 8483 6276 8576 6304
rect 7616 6264 7622 6276
rect 8570 6264 8576 6276
rect 8628 6304 8634 6316
rect 9398 6304 9404 6316
rect 8628 6276 9404 6304
rect 8628 6264 8634 6276
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12325 6307 12383 6313
rect 12325 6304 12337 6307
rect 12216 6276 12337 6304
rect 12216 6264 12222 6276
rect 12325 6273 12337 6276
rect 12371 6273 12383 6307
rect 12325 6267 12383 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 16040 6304 16068 6344
rect 14599 6276 16068 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 17034 6304 17040 6316
rect 16172 6276 16804 6304
rect 16995 6276 17040 6304
rect 16172 6264 16178 6276
rect 7098 6236 7104 6248
rect 6104 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 8389 6239 8447 6245
rect 7524 6208 7569 6236
rect 7524 6196 7530 6208
rect 8389 6205 8401 6239
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 1636 6140 2268 6168
rect 1636 6128 1642 6140
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3789 6103 3847 6109
rect 3789 6100 3801 6103
rect 3016 6072 3801 6100
rect 3016 6060 3022 6072
rect 3789 6069 3801 6072
rect 3835 6100 3847 6103
rect 4522 6100 4528 6112
rect 3835 6072 4528 6100
rect 3835 6069 3847 6072
rect 3789 6063 3847 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 5074 6100 5080 6112
rect 4663 6072 5080 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 5684 6072 6469 6100
rect 5684 6060 5690 6072
rect 6457 6069 6469 6072
rect 6503 6100 6515 6103
rect 6822 6100 6828 6112
rect 6503 6072 6828 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 8404 6100 8432 6199
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 8904 6208 9812 6236
rect 8904 6196 8910 6208
rect 8938 6168 8944 6180
rect 8899 6140 8944 6168
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9674 6168 9680 6180
rect 9232 6140 9680 6168
rect 9232 6109 9260 6140
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 8404 6072 9229 6100
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 9585 6103 9643 6109
rect 9585 6100 9597 6103
rect 9456 6072 9597 6100
rect 9456 6060 9462 6072
rect 9585 6069 9597 6072
rect 9631 6069 9643 6103
rect 9784 6100 9812 6208
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11756 6208 12081 6236
rect 11756 6196 11762 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 15746 6236 15752 6248
rect 15707 6208 15752 6236
rect 12069 6199 12127 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16390 6236 16396 6248
rect 15887 6208 16396 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16776 6245 16804 6276
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6205 16819 6239
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 16761 6199 16819 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 18156 6236 18184 6344
rect 18693 6341 18705 6375
rect 18739 6372 18751 6375
rect 19702 6372 19708 6384
rect 18739 6344 19708 6372
rect 18739 6341 18751 6344
rect 18693 6335 18751 6341
rect 19702 6332 19708 6344
rect 19760 6372 19766 6384
rect 19760 6344 20392 6372
rect 19760 6332 19766 6344
rect 20364 6316 20392 6344
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 19058 6304 19064 6316
rect 18288 6276 19064 6304
rect 18288 6264 18294 6276
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 19610 6304 19616 6316
rect 19168 6276 19616 6304
rect 18156 6208 18644 6236
rect 14921 6171 14979 6177
rect 14921 6137 14933 6171
rect 14967 6168 14979 6171
rect 17770 6168 17776 6180
rect 14967 6140 17776 6168
rect 14967 6137 14979 6140
rect 14921 6131 14979 6137
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 18230 6168 18236 6180
rect 17880 6140 18236 6168
rect 13446 6100 13452 6112
rect 9784 6072 13452 6100
rect 9585 6063 9643 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 13725 6103 13783 6109
rect 13725 6100 13737 6103
rect 13688 6072 13737 6100
rect 13688 6060 13694 6072
rect 13725 6069 13737 6072
rect 13771 6069 13783 6103
rect 13725 6063 13783 6069
rect 15289 6103 15347 6109
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 17880 6100 17908 6140
rect 18230 6128 18236 6140
rect 18288 6128 18294 6180
rect 18616 6168 18644 6208
rect 18690 6196 18696 6248
rect 18748 6236 18754 6248
rect 19168 6236 19196 6276
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 20070 6264 20076 6316
rect 20128 6313 20134 6316
rect 20128 6304 20140 6313
rect 20128 6276 20173 6304
rect 20128 6267 20140 6276
rect 20128 6264 20134 6267
rect 20346 6264 20352 6316
rect 20404 6304 20410 6316
rect 20990 6304 20996 6316
rect 20404 6276 20497 6304
rect 20951 6276 20996 6304
rect 20404 6264 20410 6276
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21358 6304 21364 6316
rect 21131 6276 21364 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 18748 6208 19196 6236
rect 18748 6196 18754 6208
rect 18966 6168 18972 6180
rect 18616 6140 18972 6168
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 21100 6168 21128 6267
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 20364 6140 21128 6168
rect 15335 6072 17908 6100
rect 17957 6103 18015 6109
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 17957 6069 17969 6103
rect 18003 6100 18015 6103
rect 18138 6100 18144 6112
rect 18003 6072 18144 6100
rect 18003 6069 18015 6072
rect 17957 6063 18015 6069
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 20364 6100 20392 6140
rect 18371 6072 20392 6100
rect 20625 6103 20683 6109
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 20625 6069 20637 6103
rect 20671 6100 20683 6103
rect 20898 6100 20904 6112
rect 20671 6072 20904 6100
rect 20671 6069 20683 6072
rect 20625 6063 20683 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 21192 6100 21220 6199
rect 21140 6072 21220 6100
rect 21140 6060 21146 6072
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4120 5868 4445 5896
rect 4120 5856 4126 5868
rect 4433 5865 4445 5868
rect 4479 5896 4491 5899
rect 4614 5896 4620 5908
rect 4479 5868 4620 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5350 5896 5356 5908
rect 5215 5868 5356 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5592 5868 5825 5896
rect 5592 5856 5598 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7432 5868 11008 5896
rect 7432 5856 7438 5868
rect 4522 5828 4528 5840
rect 3160 5800 4528 5828
rect 3160 5772 3188 5800
rect 4522 5788 4528 5800
rect 4580 5828 4586 5840
rect 5445 5831 5503 5837
rect 5445 5828 5457 5831
rect 4580 5800 5457 5828
rect 4580 5788 4586 5800
rect 5445 5797 5457 5800
rect 5491 5797 5503 5831
rect 5445 5791 5503 5797
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1728 5732 1777 5760
rect 1728 5720 1734 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 3142 5760 3148 5772
rect 3103 5732 3148 5760
rect 1765 5723 1823 5729
rect 3142 5720 3148 5732
rect 3200 5720 3206 5772
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 3970 5760 3976 5772
rect 3375 5732 3976 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 5460 5760 5488 5791
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6052 5800 9168 5828
rect 6052 5788 6058 5800
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 5460 5732 6285 5760
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 6273 5723 6331 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 7524 5732 8953 5760
rect 7524 5720 7530 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 9140 5760 9168 5800
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9585 5831 9643 5837
rect 9585 5828 9597 5831
rect 9364 5800 9597 5828
rect 9364 5788 9370 5800
rect 9585 5797 9597 5800
rect 9631 5797 9643 5831
rect 10980 5828 11008 5868
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 18598 5896 18604 5908
rect 12032 5868 18604 5896
rect 12032 5856 12038 5868
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 20346 5896 20352 5908
rect 19260 5868 20352 5896
rect 10980 5800 14596 5828
rect 9585 5791 9643 5797
rect 9140 5732 9674 5760
rect 8941 5723 8999 5729
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5442 5692 5448 5704
rect 4847 5664 5448 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5442 5652 5448 5664
rect 5500 5692 5506 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5500 5664 6193 5692
rect 5500 5652 5506 5664
rect 6181 5661 6193 5664
rect 6227 5661 6239 5695
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 6181 5655 6239 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 9646 5692 9674 5732
rect 10888 5732 11468 5760
rect 10888 5692 10916 5732
rect 9646 5664 10916 5692
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11011 5664 11376 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 2041 5627 2099 5633
rect 2041 5593 2053 5627
rect 2087 5624 2099 5627
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2087 5596 3801 5624
rect 2087 5593 2099 5596
rect 2041 5587 2099 5593
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 7558 5624 7564 5636
rect 7515 5596 7564 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 7558 5584 7564 5596
rect 7616 5624 7622 5636
rect 8389 5627 8447 5633
rect 7616 5596 7880 5624
rect 7616 5584 7622 5596
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1820 5528 1961 5556
rect 1820 5516 1826 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 1949 5519 2007 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7742 5556 7748 5568
rect 6788 5528 7748 5556
rect 6788 5516 6794 5528
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 7852 5556 7880 5596
rect 8389 5593 8401 5627
rect 8435 5624 8447 5627
rect 8662 5624 8668 5636
rect 8435 5596 8668 5624
rect 8435 5593 8447 5596
rect 8389 5587 8447 5593
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 9950 5624 9956 5636
rect 9232 5596 9956 5624
rect 9232 5556 9260 5596
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10698 5627 10756 5633
rect 10698 5624 10710 5627
rect 10100 5596 10710 5624
rect 10100 5584 10106 5596
rect 10698 5593 10710 5596
rect 10744 5593 10756 5627
rect 10698 5587 10756 5593
rect 7852 5528 9260 5556
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 10226 5556 10232 5568
rect 9364 5528 10232 5556
rect 9364 5516 9370 5528
rect 10226 5516 10232 5528
rect 10284 5556 10290 5568
rect 11238 5556 11244 5568
rect 10284 5528 11244 5556
rect 10284 5516 10290 5528
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11348 5565 11376 5664
rect 11440 5624 11468 5732
rect 13446 5720 13452 5772
rect 13504 5760 13510 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13504 5732 13645 5760
rect 13504 5720 13510 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14568 5692 14596 5800
rect 19260 5769 19288 5868
rect 20346 5856 20352 5868
rect 20404 5896 20410 5908
rect 20622 5896 20628 5908
rect 20404 5868 20628 5896
rect 20404 5856 20410 5868
rect 20622 5856 20628 5868
rect 20680 5896 20686 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20680 5868 21281 5896
rect 20680 5856 20686 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 20993 5831 21051 5837
rect 20993 5797 21005 5831
rect 21039 5828 21051 5831
rect 21174 5828 21180 5840
rect 21039 5800 21180 5828
rect 21039 5797 21051 5800
rect 20993 5791 21051 5797
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 17788 5732 18429 5760
rect 15562 5692 15568 5704
rect 14568 5664 15424 5692
rect 15523 5664 15568 5692
rect 12434 5624 12440 5636
rect 11440 5596 12440 5624
rect 12434 5584 12440 5596
rect 12492 5584 12498 5636
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 15298 5627 15356 5633
rect 15298 5624 15310 5627
rect 14516 5596 15310 5624
rect 14516 5584 14522 5596
rect 15298 5593 15310 5596
rect 15344 5593 15356 5627
rect 15396 5624 15424 5664
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5692 17558 5704
rect 17788 5701 17816 5732
rect 18417 5729 18429 5732
rect 18463 5760 18475 5763
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18463 5732 19257 5760
rect 18463 5729 18475 5732
rect 18417 5723 18475 5729
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17552 5664 17785 5692
rect 17552 5652 17558 5664
rect 17773 5661 17785 5664
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18230 5652 18236 5704
rect 18288 5692 18294 5704
rect 21008 5692 21036 5791
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 18288 5664 21036 5692
rect 18288 5652 18294 5664
rect 17218 5624 17224 5636
rect 17276 5633 17282 5636
rect 15396 5596 17224 5624
rect 15298 5587 15356 5593
rect 17218 5584 17224 5596
rect 17276 5624 17288 5633
rect 17678 5624 17684 5636
rect 17276 5596 17684 5624
rect 17276 5587 17288 5596
rect 17276 5584 17282 5587
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 19168 5596 19502 5624
rect 19168 5568 19196 5596
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 19490 5587 19548 5593
rect 11333 5559 11391 5565
rect 11333 5525 11345 5559
rect 11379 5556 11391 5559
rect 11698 5556 11704 5568
rect 11379 5528 11704 5556
rect 11379 5525 11391 5528
rect 11333 5519 11391 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13872 5528 14197 5556
rect 13872 5516 13878 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 14185 5519 14243 5525
rect 15746 5516 15752 5568
rect 15804 5556 15810 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15804 5528 16129 5556
rect 15804 5516 15810 5528
rect 16117 5525 16129 5528
rect 16163 5556 16175 5559
rect 18046 5556 18052 5568
rect 16163 5528 18052 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18877 5559 18935 5565
rect 18877 5525 18889 5559
rect 18923 5556 18935 5559
rect 19150 5556 19156 5568
rect 18923 5528 19156 5556
rect 18923 5525 18935 5528
rect 18877 5519 18935 5525
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 19702 5516 19708 5568
rect 19760 5556 19766 5568
rect 20162 5556 20168 5568
rect 19760 5528 20168 5556
rect 19760 5516 19766 5528
rect 20162 5516 20168 5528
rect 20220 5556 20226 5568
rect 20530 5556 20536 5568
rect 20220 5528 20536 5556
rect 20220 5516 20226 5528
rect 20530 5516 20536 5528
rect 20588 5556 20594 5568
rect 20625 5559 20683 5565
rect 20625 5556 20637 5559
rect 20588 5528 20637 5556
rect 20588 5516 20594 5528
rect 20625 5525 20637 5528
rect 20671 5525 20683 5559
rect 20625 5519 20683 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2590 5352 2596 5364
rect 2551 5324 2596 5352
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 3200 5324 3249 5352
rect 3200 5312 3206 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4212 5324 4261 5352
rect 4212 5312 4218 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 5258 5352 5264 5364
rect 4387 5324 5264 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 6880 5324 8861 5352
rect 6880 5312 6886 5324
rect 8849 5321 8861 5324
rect 8895 5352 8907 5355
rect 9214 5352 9220 5364
rect 8895 5324 9220 5352
rect 8895 5321 8907 5324
rect 8849 5315 8907 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 13722 5312 13728 5364
rect 13780 5312 13786 5364
rect 15286 5352 15292 5364
rect 14936 5324 15292 5352
rect 4614 5244 4620 5296
rect 4672 5284 4678 5296
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 4672 5256 5457 5284
rect 4672 5244 4678 5256
rect 5445 5253 5457 5256
rect 5491 5253 5503 5287
rect 11698 5284 11704 5296
rect 5445 5247 5503 5253
rect 9416 5256 11704 5284
rect 5353 5219 5411 5225
rect 2424 5188 3740 5216
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 2314 5148 2320 5160
rect 1627 5120 2320 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2424 5157 2452 5188
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 2516 5080 2544 5111
rect 3142 5080 3148 5092
rect 2516 5052 3148 5080
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1820 4984 1869 5012
rect 1820 4972 1826 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 2958 5012 2964 5024
rect 2919 4984 2964 5012
rect 1857 4975 1915 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3712 5021 3740 5188
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5399 5188 6377 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 7098 5216 7104 5228
rect 7059 5188 7104 5216
rect 6365 5179 6423 5185
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8386 5216 8392 5228
rect 8159 5188 8392 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 9416 5225 9444 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 13572 5287 13630 5293
rect 13572 5253 13584 5287
rect 13618 5284 13630 5287
rect 13740 5284 13768 5312
rect 13618 5256 13768 5284
rect 13618 5253 13630 5256
rect 13572 5247 13630 5253
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9668 5219 9726 5225
rect 9668 5185 9680 5219
rect 9714 5216 9726 5219
rect 10134 5216 10140 5228
rect 9714 5188 10140 5216
rect 9714 5185 9726 5188
rect 9668 5179 9726 5185
rect 10134 5176 10140 5188
rect 10192 5216 10198 5228
rect 11057 5219 11115 5225
rect 11057 5216 11069 5219
rect 10192 5188 11069 5216
rect 10192 5176 10198 5188
rect 11057 5185 11069 5188
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14936 5225 14964 5324
rect 15286 5312 15292 5324
rect 15344 5352 15350 5364
rect 15562 5352 15568 5364
rect 15344 5324 15568 5352
rect 15344 5312 15350 5324
rect 15562 5312 15568 5324
rect 15620 5352 15626 5364
rect 15657 5355 15715 5361
rect 15657 5352 15669 5355
rect 15620 5324 15669 5352
rect 15620 5312 15626 5324
rect 15657 5321 15669 5324
rect 15703 5352 15715 5355
rect 16850 5352 16856 5364
rect 15703 5324 16856 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 16850 5312 16856 5324
rect 16908 5352 16914 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16908 5324 16957 5352
rect 16908 5312 16914 5324
rect 16945 5321 16957 5324
rect 16991 5352 17003 5355
rect 17494 5352 17500 5364
rect 16991 5324 17500 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 17494 5312 17500 5324
rect 17552 5352 17558 5364
rect 17681 5355 17739 5361
rect 17681 5352 17693 5355
rect 17552 5324 17693 5352
rect 17552 5312 17558 5324
rect 17681 5321 17693 5324
rect 17727 5321 17739 5355
rect 17681 5315 17739 5321
rect 20257 5355 20315 5361
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20303 5324 21005 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 15378 5284 15384 5296
rect 15291 5256 15384 5284
rect 15378 5244 15384 5256
rect 15436 5284 15442 5296
rect 20714 5284 20720 5296
rect 15436 5256 20720 5284
rect 15436 5244 15442 5256
rect 20714 5244 20720 5256
rect 20772 5244 20778 5296
rect 20898 5284 20904 5296
rect 20859 5256 20904 5284
rect 20898 5244 20904 5256
rect 20956 5244 20962 5296
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13780 5188 13829 5216
rect 13780 5176 13786 5188
rect 13817 5185 13829 5188
rect 13863 5216 13875 5219
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13863 5188 14105 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14139 5188 14933 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 16574 5216 16580 5228
rect 14921 5179 14979 5185
rect 15672 5188 16580 5216
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4614 5148 4620 5160
rect 4203 5120 4620 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5994 5148 6000 5160
rect 5675 5120 6000 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7650 5148 7656 5160
rect 7423 5120 7656 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 15672 5148 15700 5188
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 17310 5216 17316 5228
rect 17271 5188 17316 5216
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 18966 5216 18972 5228
rect 18555 5188 18972 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 18966 5176 18972 5188
rect 19024 5216 19030 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19024 5188 19901 5216
rect 19024 5176 19030 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20530 5176 20536 5228
rect 20588 5216 20594 5228
rect 20588 5188 21128 5216
rect 20588 5176 20594 5188
rect 8297 5111 8355 5117
rect 15488 5120 15700 5148
rect 8312 5080 8340 5111
rect 11238 5080 11244 5092
rect 8312 5052 9444 5080
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3970 5012 3976 5024
rect 3743 4984 3976 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4948 4984 4997 5012
rect 4948 4972 4954 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 9416 5012 9444 5052
rect 10704 5052 11244 5080
rect 10704 5012 10732 5052
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 12492 5052 12537 5080
rect 12492 5040 12498 5052
rect 9416 4984 10732 5012
rect 4985 4975 5043 4981
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 10836 4984 10881 5012
rect 10836 4972 10842 4984
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11756 4984 11805 5012
rect 11756 4972 11762 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 14645 5015 14703 5021
rect 14645 4981 14657 5015
rect 14691 5012 14703 5015
rect 15488 5012 15516 5120
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 18230 5148 18236 5160
rect 16356 5120 18236 5148
rect 16356 5108 16362 5120
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 19150 5148 19156 5160
rect 18800 5120 19156 5148
rect 15562 5040 15568 5092
rect 15620 5080 15626 5092
rect 16209 5083 16267 5089
rect 16209 5080 16221 5083
rect 15620 5052 16221 5080
rect 15620 5040 15626 5052
rect 16209 5049 16221 5052
rect 16255 5080 16267 5083
rect 18138 5080 18144 5092
rect 16255 5052 16344 5080
rect 18051 5052 18144 5080
rect 16255 5049 16267 5052
rect 16209 5043 16267 5049
rect 14691 4984 15516 5012
rect 16316 5012 16344 5052
rect 18138 5040 18144 5052
rect 18196 5080 18202 5092
rect 18598 5080 18604 5092
rect 18196 5052 18604 5080
rect 18196 5040 18202 5052
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 18800 5012 18828 5120
rect 19150 5108 19156 5120
rect 19208 5148 19214 5160
rect 19613 5151 19671 5157
rect 19613 5148 19625 5151
rect 19208 5120 19625 5148
rect 19208 5108 19214 5120
rect 19613 5117 19625 5120
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 19797 5151 19855 5157
rect 19797 5117 19809 5151
rect 19843 5148 19855 5151
rect 20806 5148 20812 5160
rect 19843 5120 20812 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 18877 5083 18935 5089
rect 18877 5049 18889 5083
rect 18923 5080 18935 5083
rect 19058 5080 19064 5092
rect 18923 5052 19064 5080
rect 18923 5049 18935 5052
rect 18877 5043 18935 5049
rect 19058 5040 19064 5052
rect 19116 5080 19122 5092
rect 19812 5080 19840 5111
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 21100 5157 21128 5188
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 20530 5080 20536 5092
rect 19116 5052 19840 5080
rect 20491 5052 20536 5080
rect 19116 5040 19122 5052
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 19153 5015 19211 5021
rect 19153 5012 19165 5015
rect 16316 4984 19165 5012
rect 14691 4981 14703 4984
rect 14645 4975 14703 4981
rect 19153 4981 19165 4984
rect 19199 5012 19211 5015
rect 20898 5012 20904 5024
rect 19199 4984 20904 5012
rect 19199 4981 19211 4984
rect 19153 4975 19211 4981
rect 20898 4972 20904 4984
rect 20956 5012 20962 5024
rect 21082 5012 21088 5024
rect 20956 4984 21088 5012
rect 20956 4972 20962 4984
rect 21082 4972 21088 4984
rect 21140 4972 21146 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 1765 4811 1823 4817
rect 1765 4808 1777 4811
rect 1728 4780 1777 4808
rect 1728 4768 1734 4780
rect 1765 4777 1777 4780
rect 1811 4777 1823 4811
rect 2130 4808 2136 4820
rect 2091 4780 2136 4808
rect 1765 4771 1823 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2556 4780 3249 4808
rect 2556 4768 2562 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 6365 4811 6423 4817
rect 6365 4777 6377 4811
rect 6411 4808 6423 4811
rect 7098 4808 7104 4820
rect 6411 4780 7104 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9723 4780 12112 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 9766 4740 9772 4752
rect 4764 4712 5948 4740
rect 4764 4700 4770 4712
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 4062 4672 4068 4684
rect 2731 4644 4068 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4614 4672 4620 4684
rect 4575 4644 4620 4672
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5166 4672 5172 4684
rect 4847 4644 5172 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5920 4681 5948 4712
rect 6472 4712 9772 4740
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 1762 4604 1768 4616
rect 1535 4576 1768 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2464 4576 2881 4604
rect 2464 4564 2470 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 3200 4576 4261 4604
rect 3200 4564 3206 4576
rect 4249 4573 4261 4576
rect 4295 4604 4307 4607
rect 4430 4604 4436 4616
rect 4295 4576 4436 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5828 4604 5856 4635
rect 6472 4604 6500 4712
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10321 4743 10379 4749
rect 10321 4709 10333 4743
rect 10367 4740 10379 4743
rect 10410 4740 10416 4752
rect 10367 4712 10416 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 12084 4740 12112 4780
rect 12158 4768 12164 4820
rect 12216 4808 12222 4820
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 12216 4780 12265 4808
rect 12216 4768 12222 4780
rect 12253 4777 12265 4780
rect 12299 4777 12311 4811
rect 12253 4771 12311 4777
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4808 15531 4811
rect 16114 4808 16120 4820
rect 15519 4780 16120 4808
rect 15519 4777 15531 4780
rect 15473 4771 15531 4777
rect 16114 4768 16120 4780
rect 16172 4768 16178 4820
rect 17129 4811 17187 4817
rect 17129 4777 17141 4811
rect 17175 4808 17187 4811
rect 17310 4808 17316 4820
rect 17175 4780 17316 4808
rect 17175 4777 17187 4780
rect 17129 4771 17187 4777
rect 12618 4740 12624 4752
rect 12084 4712 12624 4740
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 5828 4576 6500 4604
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 6604 4576 6653 4604
rect 6604 4564 6610 4576
rect 6641 4573 6653 4576
rect 6687 4573 6699 4607
rect 8018 4604 8024 4616
rect 7979 4576 8024 4604
rect 6641 4567 6699 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 9140 4604 9168 4635
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9272 4644 9317 4672
rect 9646 4644 10057 4672
rect 9272 4632 9278 4644
rect 9646 4604 9674 4644
rect 10045 4641 10057 4644
rect 10091 4672 10103 4675
rect 10686 4672 10692 4684
rect 10091 4644 10692 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 13722 4672 13728 4684
rect 13679 4644 13728 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 13722 4632 13728 4644
rect 13780 4672 13786 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13780 4644 14105 4672
rect 13780 4632 13786 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 17144 4672 17172 4771
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 20162 4768 20168 4820
rect 20220 4808 20226 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20220 4780 20637 4808
rect 20220 4768 20226 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20898 4808 20904 4820
rect 20859 4780 20904 4808
rect 20625 4771 20683 4777
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 14093 4635 14151 4641
rect 16776 4644 17172 4672
rect 18800 4644 19257 4672
rect 11698 4604 11704 4616
rect 9140 4576 9674 4604
rect 11659 4576 11704 4604
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 16597 4607 16655 4613
rect 16597 4573 16609 4607
rect 16643 4604 16655 4607
rect 16776 4604 16804 4644
rect 16643 4576 16804 4604
rect 16643 4573 16655 4576
rect 16597 4567 16655 4573
rect 16850 4564 16856 4616
rect 16908 4604 16914 4616
rect 18800 4613 18828 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 18509 4607 18567 4613
rect 18509 4604 18521 4607
rect 16908 4576 18521 4604
rect 16908 4564 16914 4576
rect 18509 4573 18521 4576
rect 18555 4604 18567 4607
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18555 4576 18797 4604
rect 18555 4573 18567 4576
rect 18509 4567 18567 4573
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 19794 4604 19800 4616
rect 18785 4567 18843 4573
rect 18892 4576 19800 4604
rect 5997 4539 6055 4545
rect 5997 4536 6009 4539
rect 5276 4508 6009 4536
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3881 4471 3939 4477
rect 2832 4440 2877 4468
rect 2832 4428 2838 4440
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 3970 4468 3976 4480
rect 3927 4440 3976 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 3970 4428 3976 4440
rect 4028 4468 4034 4480
rect 5166 4468 5172 4480
rect 4028 4440 5172 4468
rect 4028 4428 4034 4440
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5276 4477 5304 4508
rect 5997 4505 6009 4508
rect 6043 4505 6055 4539
rect 5997 4499 6055 4505
rect 6917 4539 6975 4545
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 7190 4536 7196 4548
rect 6963 4508 7196 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 8297 4539 8355 4545
rect 8297 4505 8309 4539
rect 8343 4536 8355 4539
rect 8343 4508 10088 4536
rect 8343 4505 8355 4508
rect 8297 4499 8355 4505
rect 10060 4480 10088 4508
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 11434 4539 11492 4545
rect 11434 4536 11446 4539
rect 11204 4508 11446 4536
rect 11204 4496 11210 4508
rect 11434 4505 11446 4508
rect 11480 4505 11492 4539
rect 11434 4499 11492 4505
rect 12158 4496 12164 4548
rect 12216 4536 12222 4548
rect 13366 4539 13424 4545
rect 13366 4536 13378 4539
rect 12216 4508 13378 4536
rect 12216 4496 12222 4508
rect 13366 4505 13378 4508
rect 13412 4505 13424 4539
rect 13366 4499 13424 4505
rect 14829 4539 14887 4545
rect 14829 4505 14841 4539
rect 14875 4536 14887 4539
rect 18264 4539 18322 4545
rect 14875 4508 16528 4536
rect 14875 4505 14887 4508
rect 14829 4499 14887 4505
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 7834 4468 7840 4480
rect 7791 4440 7840 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 7834 4428 7840 4440
rect 7892 4468 7898 4480
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 7892 4440 9321 4468
rect 7892 4428 7898 4440
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 9309 4431 9367 4437
rect 10042 4428 10048 4480
rect 10100 4428 10106 4480
rect 15194 4468 15200 4480
rect 15155 4440 15200 4468
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 16500 4468 16528 4508
rect 17052 4508 18184 4536
rect 17052 4468 17080 4508
rect 16500 4440 17080 4468
rect 18156 4468 18184 4508
rect 18264 4505 18276 4539
rect 18310 4536 18322 4539
rect 18892 4536 18920 4576
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 18310 4508 18920 4536
rect 19512 4539 19570 4545
rect 18310 4505 18322 4508
rect 18264 4499 18322 4505
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 19886 4536 19892 4548
rect 19558 4508 19892 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 19886 4496 19892 4508
rect 19944 4496 19950 4548
rect 20254 4468 20260 4480
rect 18156 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 21358 4468 21364 4480
rect 21319 4440 21364 4468
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3016 4236 3801 4264
rect 3016 4224 3022 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 7926 4264 7932 4276
rect 7839 4236 7932 4264
rect 3789 4227 3847 4233
rect 7926 4224 7932 4236
rect 7984 4264 7990 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 7984 4236 8953 4264
rect 7984 4224 7990 4236
rect 8941 4233 8953 4236
rect 8987 4264 8999 4267
rect 9122 4264 9128 4276
rect 8987 4236 9128 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 10652 4236 11008 4264
rect 10652 4224 10658 4236
rect 2222 4156 2228 4208
rect 2280 4196 2286 4208
rect 3881 4199 3939 4205
rect 2280 4168 2636 4196
rect 2280 4156 2286 4168
rect 2608 4140 2636 4168
rect 3881 4165 3893 4199
rect 3927 4196 3939 4199
rect 4246 4196 4252 4208
rect 3927 4168 4252 4196
rect 3927 4165 3939 4168
rect 3881 4159 3939 4165
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 10870 4196 10876 4208
rect 10928 4205 10934 4208
rect 4672 4168 10876 4196
rect 4672 4156 4678 4168
rect 10870 4156 10876 4168
rect 10928 4159 10940 4205
rect 10980 4196 11008 4236
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 17497 4267 17555 4273
rect 15344 4236 15516 4264
rect 15344 4224 15350 4236
rect 12158 4196 12164 4208
rect 10980 4168 11836 4196
rect 10928 4156 10934 4159
rect 2498 4128 2504 4140
rect 2459 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2590 4088 2596 4140
rect 2648 4128 2654 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 2648 4100 3157 4128
rect 2648 4088 2654 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5960 4100 6377 4128
rect 5960 4088 5966 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 6604 4100 7481 4128
rect 6604 4088 6610 4100
rect 7469 4097 7481 4100
rect 7515 4128 7527 4131
rect 8478 4128 8484 4140
rect 7515 4100 8484 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 8570 4088 8576 4140
rect 8628 4128 8634 4140
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8628 4100 8861 4128
rect 8628 4088 8634 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 11149 4131 11207 4137
rect 8996 4100 11100 4128
rect 8996 4088 9002 4100
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4029 2375 4063
rect 2317 4023 2375 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2682 4060 2688 4072
rect 2455 4032 2688 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2332 3992 2360 4023
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 5810 4060 5816 4072
rect 3743 4032 5816 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3712 3992 3740 4023
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7006 4060 7012 4072
rect 6687 4032 7012 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7282 4020 7288 4072
rect 7340 4020 7346 4072
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 9582 4060 9588 4072
rect 8757 4023 8815 4029
rect 8956 4032 9588 4060
rect 2332 3964 3740 3992
rect 5994 3952 6000 4004
rect 6052 3992 6058 4004
rect 7300 3992 7328 4020
rect 6052 3964 7328 3992
rect 8297 3995 8355 4001
rect 6052 3952 6058 3964
rect 8297 3961 8309 3995
rect 8343 3992 8355 3995
rect 8772 3992 8800 4023
rect 8956 3992 8984 4032
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 11072 4060 11100 4100
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11330 4128 11336 4140
rect 11195 4100 11336 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11330 4088 11336 4100
rect 11388 4128 11394 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11388 4100 11529 4128
rect 11388 4088 11394 4100
rect 11517 4097 11529 4100
rect 11563 4128 11575 4131
rect 11698 4128 11704 4140
rect 11563 4100 11704 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11808 4128 11836 4168
rect 12084 4168 12164 4196
rect 12084 4128 12112 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 15488 4196 15516 4236
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 18138 4264 18144 4276
rect 17543 4236 18144 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 18138 4224 18144 4236
rect 18196 4264 18202 4276
rect 18598 4264 18604 4276
rect 18196 4236 18604 4264
rect 18196 4224 18202 4236
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 16209 4199 16267 4205
rect 16209 4196 16221 4199
rect 15120 4168 15424 4196
rect 15488 4168 16221 4196
rect 13078 4128 13084 4140
rect 11808 4100 12112 4128
rect 13039 4100 13084 4128
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13446 4128 13452 4140
rect 13407 4100 13452 4128
rect 13446 4088 13452 4100
rect 13504 4128 13510 4140
rect 15120 4128 15148 4168
rect 15286 4128 15292 4140
rect 15344 4137 15350 4140
rect 13504 4100 15148 4128
rect 15256 4100 15292 4128
rect 13504 4088 13510 4100
rect 15286 4088 15292 4100
rect 15344 4091 15356 4137
rect 15396 4128 15424 4168
rect 15580 4137 15608 4168
rect 16209 4165 16221 4168
rect 16255 4165 16267 4199
rect 16209 4159 16267 4165
rect 20346 4156 20352 4208
rect 20404 4156 20410 4208
rect 15565 4131 15623 4137
rect 15396 4100 15516 4128
rect 15344 4088 15350 4091
rect 15488 4060 15516 4100
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 19702 4128 19708 4140
rect 17368 4100 19708 4128
rect 17368 4088 17374 4100
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20364 4128 20392 4156
rect 20450 4131 20508 4137
rect 20450 4128 20462 4131
rect 20364 4100 20462 4128
rect 20450 4097 20462 4100
rect 20496 4097 20508 4131
rect 20450 4091 20508 4097
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 20680 4100 20729 4128
rect 20680 4088 20686 4100
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 21266 4128 21272 4140
rect 21227 4100 21272 4128
rect 20717 4091 20775 4097
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 11072 4032 14596 4060
rect 15488 4032 17601 4060
rect 9306 3992 9312 4004
rect 8343 3964 8984 3992
rect 9267 3964 9312 3992
rect 8343 3961 8355 3964
rect 8297 3955 8355 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9766 3992 9772 4004
rect 9727 3964 9772 3992
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 11977 3995 12035 4001
rect 11977 3992 11989 3995
rect 11204 3964 11989 3992
rect 11204 3952 11210 3964
rect 11977 3961 11989 3964
rect 12023 3961 12035 3995
rect 11977 3955 12035 3961
rect 1394 3924 1400 3936
rect 1355 3896 1400 3924
rect 1394 3884 1400 3896
rect 1452 3884 1458 3936
rect 1762 3924 1768 3936
rect 1723 3896 1768 3924
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 2866 3924 2872 3936
rect 2827 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4338 3924 4344 3936
rect 4295 3896 4344 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7282 3924 7288 3936
rect 7239 3896 7288 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 9398 3924 9404 3936
rect 8536 3896 9404 3924
rect 8536 3884 8542 3896
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 11164 3924 11192 3952
rect 9916 3896 11192 3924
rect 9916 3884 9922 3896
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12066 3924 12072 3936
rect 11388 3896 12072 3924
rect 11388 3884 11394 3896
rect 12066 3884 12072 3896
rect 12124 3924 12130 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12124 3896 12357 3924
rect 12124 3884 12130 3896
rect 12345 3893 12357 3896
rect 12391 3924 12403 3927
rect 13722 3924 13728 3936
rect 12391 3896 13728 3924
rect 12391 3893 12403 3896
rect 12345 3887 12403 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14185 3927 14243 3933
rect 14185 3893 14197 3927
rect 14231 3924 14243 3927
rect 14458 3924 14464 3936
rect 14231 3896 14464 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14568 3924 14596 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16206 3992 16212 4004
rect 15979 3964 16212 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 15286 3924 15292 3936
rect 14568 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3924 15350 3936
rect 15948 3924 15976 3955
rect 16206 3952 16212 3964
rect 16264 3952 16270 4004
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 16448 3964 17141 3992
rect 16448 3952 16454 3964
rect 17129 3961 17141 3964
rect 17175 3961 17187 3995
rect 17604 3992 17632 4023
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 17736 4032 17781 4060
rect 17736 4020 17742 4032
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 18969 4063 19027 4069
rect 18969 4060 18981 4063
rect 18932 4032 18981 4060
rect 18932 4020 18938 4032
rect 18969 4029 18981 4032
rect 19015 4029 19027 4063
rect 18969 4023 19027 4029
rect 18141 3995 18199 4001
rect 18141 3992 18153 3995
rect 17604 3964 18153 3992
rect 17129 3955 17187 3961
rect 18141 3961 18153 3964
rect 18187 3992 18199 3995
rect 18690 3992 18696 4004
rect 18187 3964 18696 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 18782 3952 18788 4004
rect 18840 3992 18846 4004
rect 18840 3964 19472 3992
rect 18840 3952 18846 3964
rect 15344 3896 15976 3924
rect 16853 3927 16911 3933
rect 15344 3884 15350 3896
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 17954 3924 17960 3936
rect 16899 3896 17960 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 17954 3884 17960 3896
rect 18012 3884 18018 3936
rect 19334 3924 19340 3936
rect 19295 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 19444 3924 19472 3964
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 19444 3896 21097 3924
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 2556 3692 2605 3720
rect 2556 3680 2562 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 2593 3683 2651 3689
rect 2682 3680 2688 3732
rect 2740 3720 2746 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 2740 3692 3433 3720
rect 2740 3680 2746 3692
rect 3421 3689 3433 3692
rect 3467 3720 3479 3723
rect 3970 3720 3976 3732
rect 3467 3692 3976 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 8110 3720 8116 3732
rect 5316 3692 8116 3720
rect 5316 3680 5322 3692
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 10594 3720 10600 3732
rect 8904 3692 9444 3720
rect 10555 3692 10600 3720
rect 8904 3680 8910 3692
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 1627 3624 2176 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 2148 3596 2176 3624
rect 2314 3612 2320 3664
rect 2372 3652 2378 3664
rect 5718 3652 5724 3664
rect 2372 3624 5724 3652
rect 2372 3612 2378 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 6730 3652 6736 3664
rect 6691 3624 6736 3652
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 9306 3652 9312 3664
rect 7239 3624 9312 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 9306 3612 9312 3624
rect 9364 3612 9370 3664
rect 9416 3652 9444 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 10928 3692 12265 3720
rect 10928 3680 10934 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 14366 3720 14372 3732
rect 12584 3692 14228 3720
rect 14327 3692 14372 3720
rect 12584 3680 12590 3692
rect 12066 3652 12072 3664
rect 9416 3624 10364 3652
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 2130 3584 2136 3596
rect 2091 3556 2136 3584
rect 1949 3547 2007 3553
rect 1964 3516 1992 3547
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 4338 3584 4344 3596
rect 4299 3556 4344 3584
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 5534 3584 5540 3596
rect 4571 3556 5540 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 7282 3584 7288 3596
rect 6227 3556 7288 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 10134 3584 10140 3596
rect 9631 3556 10140 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 2682 3516 2688 3528
rect 1964 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 2924 3488 4261 3516
rect 2924 3476 2930 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 4985 3519 5043 3525
rect 4985 3516 4997 3519
rect 4764 3488 4997 3516
rect 4764 3476 4770 3488
rect 4985 3485 4997 3488
rect 5031 3516 5043 3519
rect 7006 3516 7012 3528
rect 5031 3488 6408 3516
rect 6967 3488 7012 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 3050 3448 3056 3460
rect 2648 3420 3056 3448
rect 2648 3408 2654 3420
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 4798 3448 4804 3460
rect 3804 3420 4804 3448
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2271 3352 2881 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3804 3380 3832 3420
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 5902 3448 5908 3460
rect 5592 3420 5908 3448
rect 5592 3408 5598 3420
rect 5902 3408 5908 3420
rect 5960 3448 5966 3460
rect 6273 3451 6331 3457
rect 6273 3448 6285 3451
rect 5960 3420 6285 3448
rect 5960 3408 5966 3420
rect 6273 3417 6285 3420
rect 6319 3417 6331 3451
rect 6380 3448 6408 3488
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7558 3516 7564 3528
rect 7519 3488 7564 3516
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8168 3488 9352 3516
rect 8168 3476 8174 3488
rect 8846 3448 8852 3460
rect 6380 3420 8852 3448
rect 6273 3411 6331 3417
rect 8846 3408 8852 3420
rect 8904 3408 8910 3460
rect 9324 3448 9352 3488
rect 9600 3448 9628 3547
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10336 3457 10364 3624
rect 11992 3624 12072 3652
rect 11992 3593 12020 3624
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 14200 3652 14228 3692
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 16301 3723 16359 3729
rect 16301 3689 16313 3723
rect 16347 3720 16359 3723
rect 16574 3720 16580 3732
rect 16347 3692 16580 3720
rect 16347 3689 16359 3692
rect 16301 3683 16359 3689
rect 16574 3680 16580 3692
rect 16632 3720 16638 3732
rect 17586 3720 17592 3732
rect 16632 3692 17592 3720
rect 16632 3680 16638 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17862 3720 17868 3732
rect 17823 3692 17868 3720
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 20349 3723 20407 3729
rect 20349 3720 20361 3723
rect 18156 3692 20361 3720
rect 15562 3652 15568 3664
rect 14200 3624 15568 3652
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 15933 3655 15991 3661
rect 15933 3621 15945 3655
rect 15979 3652 15991 3655
rect 16666 3652 16672 3664
rect 15979 3624 16672 3652
rect 15979 3621 15991 3624
rect 15933 3615 15991 3621
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 16761 3655 16819 3661
rect 16761 3621 16773 3655
rect 16807 3652 16819 3655
rect 18046 3652 18052 3664
rect 16807 3624 18052 3652
rect 16807 3621 16819 3624
rect 16761 3615 16819 3621
rect 18046 3612 18052 3624
rect 18104 3612 18110 3664
rect 11970 3587 12028 3593
rect 11970 3553 11982 3587
rect 12016 3553 12028 3587
rect 15010 3584 15016 3596
rect 14971 3556 15016 3584
rect 11970 3547 12028 3553
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 15160 3556 15485 3584
rect 15160 3544 15166 3556
rect 15473 3553 15485 3556
rect 15519 3584 15531 3587
rect 17310 3584 17316 3596
rect 15519 3556 17172 3584
rect 17271 3556 17316 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 13633 3519 13691 3525
rect 12676 3488 13492 3516
rect 12676 3476 12682 3488
rect 9324 3420 9628 3448
rect 10321 3451 10379 3457
rect 10321 3417 10333 3451
rect 10367 3448 10379 3451
rect 11606 3448 11612 3460
rect 10367 3420 11612 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 11790 3457 11796 3460
rect 11732 3451 11796 3457
rect 11732 3417 11744 3451
rect 11778 3417 11796 3451
rect 11732 3411 11796 3417
rect 11790 3408 11796 3411
rect 11848 3408 11854 3460
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13366 3451 13424 3457
rect 13366 3448 13378 3451
rect 12492 3420 13378 3448
rect 12492 3408 12498 3420
rect 13366 3417 13378 3420
rect 13412 3417 13424 3451
rect 13464 3448 13492 3488
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13814 3516 13820 3528
rect 13679 3488 13820 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 17144 3516 17172 3556
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 17405 3587 17463 3593
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 18156 3584 18184 3692
rect 20349 3689 20361 3692
rect 20395 3689 20407 3723
rect 20349 3683 20407 3689
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18288 3624 19012 3652
rect 18288 3612 18294 3624
rect 17451 3556 18184 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 18414 3544 18420 3596
rect 18472 3584 18478 3596
rect 18800 3593 18828 3624
rect 18785 3587 18843 3593
rect 18472 3556 18644 3584
rect 18472 3544 18478 3556
rect 17862 3516 17868 3528
rect 17144 3488 17868 3516
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18616 3525 18644 3556
rect 18785 3553 18797 3587
rect 18831 3553 18843 3587
rect 18785 3547 18843 3553
rect 18874 3544 18880 3596
rect 18932 3544 18938 3596
rect 18984 3584 19012 3624
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19889 3655 19947 3661
rect 19889 3652 19901 3655
rect 19116 3624 19901 3652
rect 19116 3612 19122 3624
rect 19889 3621 19901 3624
rect 19935 3621 19947 3655
rect 19889 3615 19947 3621
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 18984 3556 19257 3584
rect 19245 3553 19257 3556
rect 19291 3553 19303 3587
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 19245 3547 19303 3553
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 18601 3519 18659 3525
rect 18012 3488 18552 3516
rect 18012 3476 18018 3488
rect 18524 3457 18552 3488
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 18892 3516 18920 3544
rect 18647 3488 18920 3516
rect 20073 3519 20131 3525
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20254 3516 20260 3528
rect 20119 3488 20260 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20714 3516 20720 3528
rect 20675 3488 20720 3516
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 21174 3516 21180 3528
rect 20855 3488 21180 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 14737 3451 14795 3457
rect 14737 3448 14749 3451
rect 13464 3420 14749 3448
rect 13366 3411 13424 3417
rect 14737 3417 14749 3420
rect 14783 3417 14795 3451
rect 14737 3411 14795 3417
rect 14829 3451 14887 3457
rect 14829 3417 14841 3451
rect 14875 3448 14887 3451
rect 18509 3451 18567 3457
rect 14875 3420 18184 3448
rect 14875 3417 14887 3420
rect 14829 3411 14887 3417
rect 3016 3352 3832 3380
rect 3881 3383 3939 3389
rect 3016 3340 3022 3352
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 3970 3380 3976 3392
rect 3927 3352 3976 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 5721 3383 5779 3389
rect 5721 3349 5733 3383
rect 5767 3380 5779 3383
rect 6365 3383 6423 3389
rect 6365 3380 6377 3383
rect 5767 3352 6377 3380
rect 5767 3349 5779 3352
rect 5721 3343 5779 3349
rect 6365 3349 6377 3352
rect 6411 3380 6423 3383
rect 6914 3380 6920 3392
rect 6411 3352 6920 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7742 3380 7748 3392
rect 7703 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8570 3380 8576 3392
rect 8531 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 8938 3380 8944 3392
rect 8899 3352 8944 3380
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 9088 3352 9321 3380
rect 9088 3340 9094 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9490 3380 9496 3392
rect 9447 3352 9496 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 16298 3340 16304 3392
rect 16356 3380 16362 3392
rect 18156 3389 18184 3420
rect 18509 3417 18521 3451
rect 18555 3417 18567 3451
rect 18509 3411 18567 3417
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 16356 3352 17509 3380
rect 16356 3340 16362 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3349 18199 3383
rect 18524 3380 18552 3411
rect 21358 3380 21364 3392
rect 18524 3352 21364 3380
rect 18141 3343 18199 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 3970 3136 3976 3188
rect 4028 3136 4034 3188
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4120 3148 4200 3176
rect 4120 3136 4126 3148
rect 2961 3111 3019 3117
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 3878 3108 3884 3120
rect 3007 3080 3884 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3040 2010 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2004 3012 2513 3040
rect 2004 3000 2010 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 2501 3003 2559 3009
rect 3712 3012 3801 3040
rect 3712 2904 3740 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 3988 3040 4016 3136
rect 4172 3108 4200 3148
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 4304 3148 4353 3176
rect 4304 3136 4310 3148
rect 4341 3145 4353 3148
rect 4387 3145 4399 3179
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4341 3139 4399 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 5960 3148 6837 3176
rect 5960 3136 5966 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 12621 3179 12679 3185
rect 7883 3148 12434 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 4709 3111 4767 3117
rect 4709 3108 4721 3111
rect 4172 3080 4721 3108
rect 4709 3077 4721 3080
rect 4755 3077 4767 3111
rect 4709 3071 4767 3077
rect 4982 3068 4988 3120
rect 5040 3068 5046 3120
rect 5629 3111 5687 3117
rect 5629 3077 5641 3111
rect 5675 3108 5687 3111
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 5675 3080 6745 3108
rect 5675 3077 5687 3080
rect 5629 3071 5687 3077
rect 6733 3077 6745 3080
rect 6779 3108 6791 3111
rect 6914 3108 6920 3120
rect 6779 3080 6920 3108
rect 6779 3077 6791 3080
rect 6733 3071 6791 3077
rect 6914 3068 6920 3080
rect 6972 3108 6978 3120
rect 8110 3108 8116 3120
rect 6972 3080 8116 3108
rect 6972 3068 6978 3080
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 9490 3068 9496 3120
rect 9548 3108 9554 3120
rect 11517 3111 11575 3117
rect 11517 3108 11529 3111
rect 9548 3080 11529 3108
rect 9548 3068 9554 3080
rect 11517 3077 11529 3080
rect 11563 3108 11575 3111
rect 12161 3111 12219 3117
rect 12161 3108 12173 3111
rect 11563 3080 12173 3108
rect 11563 3077 11575 3080
rect 11517 3071 11575 3077
rect 12161 3077 12173 3080
rect 12207 3077 12219 3111
rect 12406 3108 12434 3148
rect 12621 3145 12633 3179
rect 12667 3176 12679 3179
rect 13262 3176 13268 3188
rect 12667 3148 13124 3176
rect 13223 3148 13268 3176
rect 12667 3145 12679 3148
rect 12621 3139 12679 3145
rect 12894 3108 12900 3120
rect 12406 3080 12900 3108
rect 12161 3071 12219 3077
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 13096 3108 13124 3148
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13633 3179 13691 3185
rect 13633 3176 13645 3179
rect 13596 3148 13645 3176
rect 13596 3136 13602 3148
rect 13633 3145 13645 3148
rect 13679 3145 13691 3179
rect 16298 3176 16304 3188
rect 13633 3139 13691 3145
rect 14108 3148 16304 3176
rect 14108 3108 14136 3148
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 16669 3179 16727 3185
rect 16669 3145 16681 3179
rect 16715 3176 16727 3179
rect 16942 3176 16948 3188
rect 16715 3148 16948 3176
rect 16715 3145 16727 3148
rect 16669 3139 16727 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17083 3148 17693 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18138 3176 18144 3188
rect 18095 3148 18144 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 18966 3176 18972 3188
rect 18748 3148 18972 3176
rect 18748 3136 18754 3148
rect 18966 3136 18972 3148
rect 19024 3176 19030 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 19024 3148 19073 3176
rect 19024 3136 19030 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 19061 3139 19119 3145
rect 20622 3136 20628 3188
rect 20680 3136 20686 3188
rect 21361 3179 21419 3185
rect 21361 3145 21373 3179
rect 21407 3176 21419 3179
rect 21450 3176 21456 3188
rect 21407 3148 21456 3176
rect 21407 3145 21419 3148
rect 21361 3139 21419 3145
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 13096 3080 14136 3108
rect 14185 3111 14243 3117
rect 14185 3077 14197 3111
rect 14231 3108 14243 3111
rect 14231 3080 15608 3108
rect 14231 3077 14243 3080
rect 14185 3071 14243 3077
rect 4065 3043 4123 3049
rect 4065 3040 4077 3043
rect 3988 3012 4077 3040
rect 3789 3003 3847 3009
rect 4065 3009 4077 3012
rect 4111 3009 4123 3043
rect 5000 3040 5028 3068
rect 7650 3040 7656 3052
rect 5000 3012 5304 3040
rect 7611 3012 7656 3040
rect 4065 3003 4123 3009
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5166 2972 5172 2984
rect 5031 2944 5172 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5276 2972 5304 3012
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 8202 3040 8208 3052
rect 8163 3012 8208 3040
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10882 3043 10940 3049
rect 10882 3040 10894 3043
rect 9824 3012 10894 3040
rect 9824 3000 9830 3012
rect 10882 3009 10894 3012
rect 10928 3009 10940 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 10882 3003 10940 3009
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11756 3012 12265 3040
rect 11756 3000 11762 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 13909 3043 13967 3049
rect 12253 3003 12311 3009
rect 13004 3012 13308 3040
rect 7009 2975 7067 2981
rect 5276 2944 6408 2972
rect 5626 2904 5632 2916
rect 3712 2876 5632 2904
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 6380 2913 6408 2944
rect 7009 2941 7021 2975
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 10134 2972 10140 2984
rect 9079 2944 10140 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 6365 2907 6423 2913
rect 6365 2873 6377 2907
rect 6411 2873 6423 2907
rect 7024 2904 7052 2935
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12434 2972 12440 2984
rect 12069 2935 12127 2941
rect 12268 2944 12440 2972
rect 8389 2907 8447 2913
rect 7024 2876 7144 2904
rect 6365 2867 6423 2873
rect 2130 2836 2136 2848
rect 2091 2808 2136 2836
rect 2130 2796 2136 2808
rect 2188 2796 2194 2848
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 3237 2839 3295 2845
rect 3237 2836 3249 2839
rect 3016 2808 3249 2836
rect 3016 2796 3022 2808
rect 3237 2805 3249 2808
rect 3283 2805 3295 2839
rect 3237 2799 3295 2805
rect 3326 2796 3332 2848
rect 3384 2836 3390 2848
rect 5350 2836 5356 2848
rect 3384 2808 5356 2836
rect 3384 2796 3390 2808
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5776 2808 6009 2836
rect 5776 2796 5782 2808
rect 5997 2805 6009 2808
rect 6043 2836 6055 2839
rect 7116 2836 7144 2876
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 12084 2904 12112 2935
rect 12268 2904 12296 2944
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 13004 2981 13032 3012
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2941 13047 2975
rect 13170 2972 13176 2984
rect 13131 2944 13176 2972
rect 12989 2935 13047 2941
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 13280 2972 13308 3012
rect 13909 3009 13921 3043
rect 13955 3040 13967 3043
rect 14274 3040 14280 3052
rect 13955 3012 14280 3040
rect 13955 3009 13967 3012
rect 13909 3003 13967 3009
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15580 3049 15608 3080
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 16022 3108 16028 3120
rect 15804 3080 16028 3108
rect 15804 3068 15810 3080
rect 16022 3068 16028 3080
rect 16080 3108 16086 3120
rect 16117 3111 16175 3117
rect 16117 3108 16129 3111
rect 16080 3080 16129 3108
rect 16080 3068 16086 3080
rect 16117 3077 16129 3080
rect 16163 3077 16175 3111
rect 18598 3108 18604 3120
rect 16117 3071 16175 3077
rect 16500 3080 18604 3108
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14792 3012 14841 3040
rect 14792 3000 14798 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 14182 2972 14188 2984
rect 13280 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15194 2932 15200 2984
rect 15252 2972 15258 2984
rect 16500 2972 16528 3080
rect 18598 3068 18604 3080
rect 18656 3108 18662 3120
rect 19153 3111 19211 3117
rect 19153 3108 19165 3111
rect 18656 3080 19165 3108
rect 18656 3068 18662 3080
rect 19153 3077 19165 3080
rect 19199 3077 19211 3111
rect 20640 3108 20668 3136
rect 20809 3111 20867 3117
rect 20809 3108 20821 3111
rect 20640 3080 20821 3108
rect 19153 3071 19211 3077
rect 20809 3077 20821 3080
rect 20855 3077 20867 3111
rect 20809 3071 20867 3077
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 18012 3012 18153 3040
rect 18012 3000 18018 3012
rect 18141 3009 18153 3012
rect 18187 3040 18199 3043
rect 18874 3040 18880 3052
rect 18187 3012 18880 3040
rect 18187 3009 18199 3012
rect 18141 3003 18199 3009
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19978 3040 19984 3052
rect 19939 3012 19984 3040
rect 19978 3000 19984 3012
rect 20036 3040 20042 3052
rect 20622 3040 20628 3052
rect 20036 3012 20628 3040
rect 20036 3000 20042 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 15252 2944 16528 2972
rect 17129 2975 17187 2981
rect 15252 2932 15258 2944
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 14734 2904 14740 2916
rect 8435 2876 10272 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 9674 2836 9680 2848
rect 6043 2808 9680 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 10244 2836 10272 2876
rect 11164 2876 12020 2904
rect 12084 2876 12296 2904
rect 12406 2876 14740 2904
rect 11164 2836 11192 2876
rect 9824 2808 9869 2836
rect 10244 2808 11192 2836
rect 11992 2836 12020 2876
rect 12406 2836 12434 2876
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 15654 2864 15660 2916
rect 15712 2864 15718 2916
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2904 15807 2907
rect 16206 2904 16212 2916
rect 15795 2876 16212 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 17144 2904 17172 2935
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 18325 2975 18383 2981
rect 17276 2944 17321 2972
rect 17276 2932 17282 2944
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 19245 2975 19303 2981
rect 18371 2944 18920 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 18693 2907 18751 2913
rect 18693 2904 18705 2907
rect 17144 2876 18705 2904
rect 18693 2873 18705 2876
rect 18739 2873 18751 2907
rect 18892 2904 18920 2944
rect 19245 2941 19257 2975
rect 19291 2972 19303 2975
rect 19794 2972 19800 2984
rect 19291 2944 19800 2972
rect 19291 2941 19303 2944
rect 19245 2935 19303 2941
rect 19260 2904 19288 2935
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 18892 2876 19288 2904
rect 18693 2867 18751 2873
rect 11992 2808 12434 2836
rect 9824 2796 9830 2808
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 15672 2836 15700 2864
rect 14332 2808 15700 2836
rect 14332 2796 14338 2808
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 2832 2604 4077 2632
rect 2832 2592 2838 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 4065 2595 4123 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 11146 2632 11152 2644
rect 9815 2604 11152 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12529 2635 12587 2641
rect 12529 2632 12541 2635
rect 12492 2604 12541 2632
rect 12492 2592 12498 2604
rect 12529 2601 12541 2604
rect 12575 2601 12587 2635
rect 12529 2595 12587 2601
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 13170 2632 13176 2644
rect 12943 2604 13176 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 14274 2632 14280 2644
rect 14231 2604 14280 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 15194 2632 15200 2644
rect 14599 2604 15200 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 2130 2524 2136 2576
rect 2188 2564 2194 2576
rect 13262 2564 13268 2576
rect 2188 2536 13268 2564
rect 2188 2524 2194 2536
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 14568 2564 14596 2595
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17218 2592 17224 2644
rect 17276 2632 17282 2644
rect 18509 2635 18567 2641
rect 18509 2632 18521 2635
rect 17276 2604 18521 2632
rect 17276 2592 17282 2604
rect 18509 2601 18521 2604
rect 18555 2601 18567 2635
rect 18509 2595 18567 2601
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20625 2635 20683 2641
rect 20625 2632 20637 2635
rect 20496 2604 20637 2632
rect 20496 2592 20502 2604
rect 20625 2601 20637 2604
rect 20671 2601 20683 2635
rect 20625 2595 20683 2601
rect 13372 2536 14596 2564
rect 1670 2456 1676 2508
rect 1728 2496 1734 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 1728 2468 4629 2496
rect 1728 2456 1734 2468
rect 4617 2465 4629 2468
rect 4663 2496 4675 2499
rect 5258 2496 5264 2508
rect 4663 2468 5264 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 5258 2456 5264 2468
rect 5316 2496 5322 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5316 2468 5641 2496
rect 5316 2456 5322 2468
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7558 2496 7564 2508
rect 6779 2468 7564 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 12158 2496 12164 2508
rect 8628 2468 12164 2496
rect 8628 2456 8634 2468
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 13372 2505 13400 2536
rect 18414 2524 18420 2576
rect 18472 2564 18478 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 18472 2536 19349 2564
rect 18472 2524 18478 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2465 13415 2499
rect 13357 2459 13415 2465
rect 13538 2456 13544 2508
rect 13596 2496 13602 2508
rect 15654 2496 15660 2508
rect 13596 2468 15660 2496
rect 13596 2456 13602 2468
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 21174 2496 21180 2508
rect 16991 2468 17448 2496
rect 21135 2468 21180 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5592 2400 5917 2428
rect 5592 2388 5598 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 6914 2428 6920 2440
rect 6875 2400 6920 2428
rect 5905 2391 5963 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 4706 2360 4712 2372
rect 4571 2332 4712 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4706 2320 4712 2332
rect 4764 2320 4770 2372
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 7852 2360 7880 2391
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8720 2400 8953 2428
rect 8720 2388 8726 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10192 2400 10701 2428
rect 10192 2388 10198 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11296 2400 11713 2428
rect 11296 2388 11302 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 14366 2428 14372 2440
rect 11701 2391 11759 2397
rect 12406 2400 14372 2428
rect 9140 2360 9168 2388
rect 9490 2360 9496 2372
rect 5684 2332 7880 2360
rect 8864 2332 9496 2360
rect 5684 2320 5690 2332
rect 8864 2304 8892 2332
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 12406 2360 12434 2400
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 15102 2428 15108 2440
rect 15063 2400 15108 2428
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2428 15807 2431
rect 15838 2428 15844 2440
rect 15795 2400 15844 2428
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17420 2437 17448 2468
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 17405 2431 17463 2437
rect 17405 2397 17417 2431
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18322 2428 18328 2440
rect 18279 2400 18328 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 18932 2400 19533 2428
rect 18932 2388 18938 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20162 2428 20168 2440
rect 20119 2400 20168 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 20990 2428 20996 2440
rect 20951 2400 20996 2428
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 10244 2332 12434 2360
rect 13265 2363 13323 2369
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2292 3482 2304
rect 4433 2295 4491 2301
rect 4433 2292 4445 2295
rect 3476 2264 4445 2292
rect 3476 2252 3482 2264
rect 4433 2261 4445 2264
rect 4479 2261 4491 2295
rect 4433 2255 4491 2261
rect 7377 2295 7435 2301
rect 7377 2261 7389 2295
rect 7423 2292 7435 2295
rect 7834 2292 7840 2304
rect 7423 2264 7840 2292
rect 7423 2261 7435 2264
rect 7377 2255 7435 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 8018 2292 8024 2304
rect 7979 2264 8024 2292
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 8573 2295 8631 2301
rect 8573 2261 8585 2295
rect 8619 2292 8631 2295
rect 8846 2292 8852 2304
rect 8619 2264 8852 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 10134 2292 10140 2304
rect 9171 2264 10140 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 10244 2301 10272 2332
rect 13265 2329 13277 2363
rect 13311 2360 13323 2363
rect 15010 2360 15016 2372
rect 13311 2332 15016 2360
rect 13311 2329 13323 2332
rect 13265 2323 13323 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 16942 2360 16948 2372
rect 15304 2332 16948 2360
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2261 10287 2295
rect 10870 2292 10876 2304
rect 10831 2264 10876 2292
rect 10229 2255 10287 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 15194 2292 15200 2304
rect 11931 2264 15200 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 15304 2301 15332 2332
rect 16942 2320 16948 2332
rect 17000 2320 17006 2372
rect 18598 2320 18604 2372
rect 18656 2360 18662 2372
rect 18656 2332 21128 2360
rect 18656 2320 18662 2332
rect 21100 2304 21128 2332
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15933 2295 15991 2301
rect 15933 2261 15945 2295
rect 15979 2292 15991 2295
rect 16390 2292 16396 2304
rect 15979 2264 16396 2292
rect 15979 2261 15991 2264
rect 15933 2255 15991 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17368 2264 17601 2292
rect 17368 2252 17374 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17736 2264 18061 2292
rect 17736 2252 17742 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 20254 2292 20260 2304
rect 20215 2264 20260 2292
rect 18049 2255 18107 2261
rect 20254 2252 20260 2264
rect 20312 2252 20318 2304
rect 21082 2292 21088 2304
rect 21043 2264 21088 2292
rect 21082 2252 21088 2264
rect 21140 2252 21146 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 8018 2048 8024 2100
rect 8076 2088 8082 2100
rect 12526 2088 12532 2100
rect 8076 2060 12532 2088
rect 8076 2048 8082 2060
rect 12526 2048 12532 2060
rect 12584 2048 12590 2100
rect 13262 2048 13268 2100
rect 13320 2088 13326 2100
rect 19518 2088 19524 2100
rect 13320 2060 19524 2088
rect 13320 2048 13326 2060
rect 19518 2048 19524 2060
rect 19576 2048 19582 2100
rect 10870 1980 10876 2032
rect 10928 2020 10934 2032
rect 15838 2020 15844 2032
rect 10928 1992 15844 2020
rect 10928 1980 10934 1992
rect 15838 1980 15844 1992
rect 15896 1980 15902 2032
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 13262 1952 13268 1964
rect 7892 1924 13268 1952
rect 7892 1912 7898 1924
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 10134 1844 10140 1896
rect 10192 1884 10198 1896
rect 15102 1884 15108 1896
rect 10192 1856 15108 1884
rect 10192 1844 10198 1856
rect 15102 1844 15108 1856
rect 15160 1844 15166 1896
rect 7282 1776 7288 1828
rect 7340 1816 7346 1828
rect 13538 1816 13544 1828
rect 7340 1788 13544 1816
rect 7340 1776 7346 1788
rect 13538 1776 13544 1788
rect 13596 1776 13602 1828
rect 9582 1640 9588 1692
rect 9640 1680 9646 1692
rect 10502 1680 10508 1692
rect 9640 1652 10508 1680
rect 9640 1640 9646 1652
rect 10502 1640 10508 1652
rect 10560 1640 10566 1692
rect 9306 1368 9312 1420
rect 9364 1408 9370 1420
rect 13630 1408 13636 1420
rect 9364 1380 13636 1408
rect 9364 1368 9370 1380
rect 13630 1368 13636 1380
rect 13688 1368 13694 1420
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 20260 20544 20312 20596
rect 13728 20476 13780 20528
rect 14372 20408 14424 20460
rect 7840 20383 7892 20392
rect 7840 20349 7849 20383
rect 7849 20349 7883 20383
rect 7883 20349 7892 20383
rect 7840 20340 7892 20349
rect 18236 20408 18288 20460
rect 19892 20408 19944 20460
rect 18144 20340 18196 20392
rect 4068 20204 4120 20256
rect 12348 20247 12400 20256
rect 12348 20213 12357 20247
rect 12357 20213 12391 20247
rect 12391 20213 12400 20247
rect 12348 20204 12400 20213
rect 17408 20247 17460 20256
rect 17408 20213 17417 20247
rect 17417 20213 17451 20247
rect 17451 20213 17460 20247
rect 17408 20204 17460 20213
rect 18144 20204 18196 20256
rect 18512 20204 18564 20256
rect 19892 20247 19944 20256
rect 19892 20213 19901 20247
rect 19901 20213 19935 20247
rect 19935 20213 19944 20247
rect 19892 20204 19944 20213
rect 20444 20247 20496 20256
rect 20444 20213 20453 20247
rect 20453 20213 20487 20247
rect 20487 20213 20496 20247
rect 20444 20204 20496 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2780 20000 2832 20052
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 14372 20000 14424 20052
rect 14556 20000 14608 20052
rect 18052 20000 18104 20052
rect 20628 20000 20680 20052
rect 8484 19864 8536 19916
rect 10508 19907 10560 19916
rect 10508 19873 10517 19907
rect 10517 19873 10551 19907
rect 10551 19873 10560 19907
rect 10508 19864 10560 19873
rect 3884 19796 3936 19848
rect 4712 19796 4764 19848
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 9864 19796 9916 19848
rect 11060 19796 11112 19848
rect 12624 19932 12676 19984
rect 17960 19932 18012 19984
rect 12440 19864 12492 19916
rect 12348 19796 12400 19848
rect 13728 19864 13780 19916
rect 14740 19907 14792 19916
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 16028 19864 16080 19916
rect 17684 19864 17736 19916
rect 18236 19907 18288 19916
rect 18236 19873 18245 19907
rect 18245 19873 18279 19907
rect 18279 19873 18288 19907
rect 18236 19864 18288 19873
rect 13636 19796 13688 19848
rect 14832 19796 14884 19848
rect 17408 19796 17460 19848
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 7932 19660 7984 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 11060 19703 11112 19712
rect 10416 19660 10468 19669
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11888 19728 11940 19780
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 14556 19660 14608 19712
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 16948 19660 17000 19712
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 17592 19660 17644 19669
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2872 19456 2924 19508
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 7932 19499 7984 19508
rect 7932 19465 7941 19499
rect 7941 19465 7975 19499
rect 7975 19465 7984 19499
rect 7932 19456 7984 19465
rect 10416 19499 10468 19508
rect 10416 19465 10425 19499
rect 10425 19465 10459 19499
rect 10459 19465 10468 19499
rect 10416 19456 10468 19465
rect 11704 19456 11756 19508
rect 12624 19456 12676 19508
rect 14832 19499 14884 19508
rect 14372 19431 14424 19440
rect 14372 19397 14381 19431
rect 14381 19397 14415 19431
rect 14415 19397 14424 19431
rect 14372 19388 14424 19397
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 16028 19499 16080 19508
rect 16028 19465 16037 19499
rect 16037 19465 16071 19499
rect 16071 19465 16080 19499
rect 16028 19456 16080 19465
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 17592 19456 17644 19508
rect 18696 19456 18748 19508
rect 18512 19388 18564 19440
rect 2504 19320 2556 19372
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 5172 19363 5224 19372
rect 5172 19329 5181 19363
rect 5181 19329 5215 19363
rect 5215 19329 5224 19363
rect 5172 19320 5224 19329
rect 8576 19320 8628 19372
rect 3976 19252 4028 19304
rect 1952 19227 2004 19236
rect 1952 19193 1961 19227
rect 1961 19193 1995 19227
rect 1995 19193 2004 19227
rect 1952 19184 2004 19193
rect 7288 19252 7340 19304
rect 8024 19295 8076 19304
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 9312 19252 9364 19304
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 15384 19320 15436 19372
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 10140 19252 10192 19304
rect 12348 19295 12400 19304
rect 12348 19261 12357 19295
rect 12357 19261 12391 19295
rect 12391 19261 12400 19295
rect 12348 19252 12400 19261
rect 15476 19252 15528 19304
rect 6552 19116 6604 19168
rect 7564 19159 7616 19168
rect 7564 19125 7573 19159
rect 7573 19125 7607 19159
rect 7607 19125 7616 19159
rect 7564 19116 7616 19125
rect 15200 19116 15252 19168
rect 16488 19184 16540 19236
rect 17776 19252 17828 19304
rect 17224 19116 17276 19168
rect 17868 19116 17920 19168
rect 20904 19159 20956 19168
rect 20904 19125 20913 19159
rect 20913 19125 20947 19159
rect 20947 19125 20956 19159
rect 20904 19116 20956 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 5080 18912 5132 18964
rect 5080 18776 5132 18828
rect 6552 18776 6604 18828
rect 6828 18776 6880 18828
rect 8944 18819 8996 18828
rect 8944 18785 8953 18819
rect 8953 18785 8987 18819
rect 8987 18785 8996 18819
rect 13544 18912 13596 18964
rect 14464 18912 14516 18964
rect 14648 18912 14700 18964
rect 16488 18912 16540 18964
rect 16948 18912 17000 18964
rect 17776 18912 17828 18964
rect 18328 18912 18380 18964
rect 18512 18955 18564 18964
rect 18512 18921 18521 18955
rect 18521 18921 18555 18955
rect 18555 18921 18564 18955
rect 18512 18912 18564 18921
rect 12072 18844 12124 18896
rect 12440 18844 12492 18896
rect 8944 18776 8996 18785
rect 10968 18776 11020 18828
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 18696 18844 18748 18896
rect 20812 18844 20864 18896
rect 4252 18708 4304 18760
rect 1768 18640 1820 18692
rect 8300 18708 8352 18760
rect 11612 18708 11664 18760
rect 12348 18708 12400 18760
rect 16120 18819 16172 18828
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 3148 18572 3200 18624
rect 4528 18572 4580 18624
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 5908 18572 5960 18624
rect 7288 18640 7340 18692
rect 10324 18640 10376 18692
rect 6552 18572 6604 18624
rect 7196 18572 7248 18624
rect 9680 18572 9732 18624
rect 9956 18572 10008 18624
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 11244 18572 11296 18624
rect 11704 18640 11756 18692
rect 12072 18572 12124 18624
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 15016 18708 15068 18760
rect 16120 18785 16129 18819
rect 16129 18785 16163 18819
rect 16163 18785 16172 18819
rect 16120 18776 16172 18785
rect 17132 18776 17184 18828
rect 18144 18776 18196 18828
rect 15200 18708 15252 18760
rect 16212 18708 16264 18760
rect 18236 18708 18288 18760
rect 18604 18708 18656 18760
rect 20168 18776 20220 18828
rect 19800 18708 19852 18760
rect 16396 18640 16448 18692
rect 16948 18683 17000 18692
rect 16948 18649 16957 18683
rect 16957 18649 16991 18683
rect 16991 18649 17000 18683
rect 16948 18640 17000 18649
rect 18052 18683 18104 18692
rect 18052 18649 18061 18683
rect 18061 18649 18095 18683
rect 18095 18649 18104 18683
rect 18052 18640 18104 18649
rect 18880 18640 18932 18692
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 15384 18572 15436 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 17500 18572 17552 18624
rect 19432 18572 19484 18624
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 19616 18572 19668 18581
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 7288 18368 7340 18420
rect 8024 18368 8076 18420
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 8484 18368 8536 18420
rect 10048 18368 10100 18420
rect 6920 18300 6972 18352
rect 12808 18368 12860 18420
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 4068 18232 4120 18284
rect 6000 18232 6052 18284
rect 8668 18232 8720 18284
rect 8944 18232 8996 18284
rect 3148 18207 3200 18216
rect 1584 18028 1636 18080
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 3148 18173 3157 18207
rect 3157 18173 3191 18207
rect 3191 18173 3200 18207
rect 3148 18164 3200 18173
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 4804 18164 4856 18216
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 8484 18207 8536 18216
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 8484 18164 8536 18173
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 17408 18300 17460 18352
rect 17500 18300 17552 18352
rect 18512 18368 18564 18420
rect 19156 18343 19208 18352
rect 19156 18309 19165 18343
rect 19165 18309 19199 18343
rect 19199 18309 19208 18343
rect 19156 18300 19208 18309
rect 19432 18300 19484 18352
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 13544 18232 13596 18284
rect 13728 18232 13780 18284
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 18328 18232 18380 18284
rect 20352 18232 20404 18284
rect 21272 18232 21324 18284
rect 9496 18164 9548 18173
rect 11888 18207 11940 18216
rect 4344 18096 4396 18148
rect 5816 18096 5868 18148
rect 8300 18096 8352 18148
rect 11888 18173 11897 18207
rect 11897 18173 11931 18207
rect 11931 18173 11940 18207
rect 11888 18164 11940 18173
rect 14464 18164 14516 18216
rect 17408 18164 17460 18216
rect 16948 18096 17000 18148
rect 4436 18028 4488 18080
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 6644 18071 6696 18080
rect 6644 18037 6653 18071
rect 6653 18037 6687 18071
rect 6687 18037 6696 18071
rect 6644 18028 6696 18037
rect 7380 18028 7432 18080
rect 8484 18028 8536 18080
rect 10324 18028 10376 18080
rect 10784 18028 10836 18080
rect 14740 18028 14792 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 16304 18028 16356 18080
rect 18236 18028 18288 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 19064 18164 19116 18216
rect 18972 18096 19024 18148
rect 19432 18028 19484 18080
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 20444 18028 20496 18037
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1860 17824 1912 17876
rect 2780 17824 2832 17876
rect 5172 17824 5224 17876
rect 6000 17824 6052 17876
rect 8760 17824 8812 17876
rect 9404 17824 9456 17876
rect 9772 17824 9824 17876
rect 15200 17824 15252 17876
rect 16488 17824 16540 17876
rect 17776 17824 17828 17876
rect 19064 17824 19116 17876
rect 19340 17824 19392 17876
rect 21272 17867 21324 17876
rect 3240 17688 3292 17740
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 11060 17756 11112 17808
rect 12348 17756 12400 17808
rect 16396 17756 16448 17808
rect 4804 17688 4856 17697
rect 6920 17731 6972 17740
rect 2412 17620 2464 17672
rect 6920 17697 6929 17731
rect 6929 17697 6963 17731
rect 6963 17697 6972 17731
rect 6920 17688 6972 17697
rect 9496 17688 9548 17740
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 10692 17688 10744 17740
rect 18236 17731 18288 17740
rect 18236 17697 18245 17731
rect 18245 17697 18279 17731
rect 18279 17697 18288 17731
rect 18236 17688 18288 17697
rect 18420 17688 18472 17740
rect 6552 17620 6604 17672
rect 15844 17620 15896 17672
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 18052 17620 18104 17672
rect 19892 17688 19944 17740
rect 21272 17833 21281 17867
rect 21281 17833 21315 17867
rect 21315 17833 21324 17867
rect 21272 17824 21324 17833
rect 4804 17552 4856 17604
rect 5724 17552 5776 17604
rect 7380 17552 7432 17604
rect 9404 17552 9456 17604
rect 9772 17552 9824 17604
rect 10324 17552 10376 17604
rect 10600 17552 10652 17604
rect 14280 17552 14332 17604
rect 20720 17620 20772 17672
rect 1676 17484 1728 17536
rect 2964 17484 3016 17536
rect 4988 17527 5040 17536
rect 4988 17493 4997 17527
rect 4997 17493 5031 17527
rect 5031 17493 5040 17527
rect 4988 17484 5040 17493
rect 5172 17484 5224 17536
rect 6000 17527 6052 17536
rect 6000 17493 6009 17527
rect 6009 17493 6043 17527
rect 6043 17493 6052 17527
rect 6000 17484 6052 17493
rect 6552 17484 6604 17536
rect 6644 17484 6696 17536
rect 7012 17527 7064 17536
rect 7012 17493 7021 17527
rect 7021 17493 7055 17527
rect 7055 17493 7064 17527
rect 7012 17484 7064 17493
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7472 17527 7524 17536
rect 7104 17484 7156 17493
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 8392 17484 8444 17536
rect 8760 17484 8812 17536
rect 9588 17484 9640 17536
rect 9680 17484 9732 17536
rect 10416 17484 10468 17536
rect 13544 17484 13596 17536
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 19984 17484 20036 17536
rect 20444 17484 20496 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 20904 17484 20956 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1492 17323 1544 17332
rect 1492 17289 1501 17323
rect 1501 17289 1535 17323
rect 1535 17289 1544 17323
rect 1492 17280 1544 17289
rect 3884 17280 3936 17332
rect 4068 17280 4120 17332
rect 4160 17280 4212 17332
rect 5172 17323 5224 17332
rect 5172 17289 5181 17323
rect 5181 17289 5215 17323
rect 5215 17289 5224 17323
rect 5172 17280 5224 17289
rect 5816 17280 5868 17332
rect 8392 17323 8444 17332
rect 3332 17212 3384 17264
rect 4620 17212 4672 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 1584 17008 1636 17060
rect 4436 17076 4488 17128
rect 2136 16983 2188 16992
rect 2136 16949 2145 16983
rect 2145 16949 2179 16983
rect 2179 16949 2188 16983
rect 2136 16940 2188 16949
rect 2872 16940 2924 16992
rect 3056 16940 3108 16992
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 8392 17289 8401 17323
rect 8401 17289 8435 17323
rect 8435 17289 8444 17323
rect 8392 17280 8444 17289
rect 8484 17323 8536 17332
rect 8484 17289 8493 17323
rect 8493 17289 8527 17323
rect 8527 17289 8536 17323
rect 8484 17280 8536 17289
rect 8668 17280 8720 17332
rect 9956 17280 10008 17332
rect 10416 17280 10468 17332
rect 10600 17280 10652 17332
rect 14280 17323 14332 17332
rect 9588 17212 9640 17264
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 8668 17119 8720 17128
rect 7840 17008 7892 17060
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 5816 16940 5868 16992
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 8392 17008 8444 17060
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 14280 17289 14289 17323
rect 14289 17289 14323 17323
rect 14323 17289 14332 17323
rect 14280 17280 14332 17289
rect 15292 17280 15344 17332
rect 15844 17280 15896 17332
rect 16856 17280 16908 17332
rect 18696 17280 18748 17332
rect 20812 17323 20864 17332
rect 13820 17212 13872 17264
rect 18052 17212 18104 17264
rect 19800 17255 19852 17264
rect 19800 17221 19809 17255
rect 19809 17221 19843 17255
rect 19843 17221 19852 17255
rect 19800 17212 19852 17221
rect 20812 17289 20821 17323
rect 20821 17289 20855 17323
rect 20855 17289 20864 17323
rect 20812 17280 20864 17289
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 16948 17144 17000 17196
rect 20076 17187 20128 17196
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 20812 17076 20864 17128
rect 15384 17008 15436 17060
rect 16120 17008 16172 17060
rect 17960 17008 18012 17060
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 12992 16940 13044 16992
rect 13268 16940 13320 16992
rect 14280 16940 14332 16992
rect 16948 16940 17000 16992
rect 18604 16940 18656 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1676 16736 1728 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 3884 16736 3936 16788
rect 5816 16736 5868 16788
rect 6920 16736 6972 16788
rect 7196 16779 7248 16788
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 8392 16736 8444 16788
rect 4528 16711 4580 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 4160 16600 4212 16652
rect 4528 16677 4537 16711
rect 4537 16677 4571 16711
rect 4571 16677 4580 16711
rect 4528 16668 4580 16677
rect 5448 16668 5500 16720
rect 7104 16668 7156 16720
rect 8300 16668 8352 16720
rect 8760 16668 8812 16720
rect 9404 16668 9456 16720
rect 2044 16464 2096 16516
rect 4712 16532 4764 16584
rect 7012 16600 7064 16652
rect 7380 16600 7432 16652
rect 7932 16600 7984 16652
rect 3424 16464 3476 16516
rect 4344 16464 4396 16516
rect 5356 16464 5408 16516
rect 5816 16507 5868 16516
rect 5816 16473 5825 16507
rect 5825 16473 5859 16507
rect 5859 16473 5868 16507
rect 5816 16464 5868 16473
rect 6644 16464 6696 16516
rect 6920 16532 6972 16584
rect 10968 16600 11020 16652
rect 15660 16736 15712 16788
rect 15752 16736 15804 16788
rect 20076 16736 20128 16788
rect 11152 16668 11204 16720
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 21088 16668 21140 16720
rect 15476 16600 15528 16652
rect 16396 16600 16448 16652
rect 16948 16600 17000 16652
rect 17040 16600 17092 16652
rect 20444 16643 20496 16652
rect 20444 16609 20453 16643
rect 20453 16609 20487 16643
rect 20487 16609 20496 16643
rect 20444 16600 20496 16609
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 18604 16532 18656 16584
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 20628 16532 20680 16584
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 4896 16396 4948 16405
rect 5080 16396 5132 16448
rect 5724 16396 5776 16448
rect 6828 16396 6880 16448
rect 7104 16464 7156 16516
rect 7012 16396 7064 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 15568 16464 15620 16516
rect 16028 16464 16080 16516
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 16396 16396 16448 16448
rect 17960 16464 18012 16516
rect 20720 16464 20772 16516
rect 18052 16396 18104 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2780 16192 2832 16244
rect 4988 16192 5040 16244
rect 5816 16192 5868 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 6828 16192 6880 16244
rect 7656 16192 7708 16244
rect 3976 16124 4028 16176
rect 7012 16167 7064 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4620 16056 4672 16108
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 4896 15988 4948 16040
rect 5264 15988 5316 16040
rect 5448 16056 5500 16108
rect 5816 15920 5868 15972
rect 1400 15852 1452 15904
rect 4344 15852 4396 15904
rect 7012 16133 7021 16167
rect 7021 16133 7055 16167
rect 7055 16133 7064 16167
rect 7012 16124 7064 16133
rect 8116 16124 8168 16176
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7380 16056 7432 16108
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 8024 16031 8076 16040
rect 7104 15988 7156 15997
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 9772 16192 9824 16244
rect 10140 16192 10192 16244
rect 12072 16192 12124 16244
rect 13452 16192 13504 16244
rect 13728 16192 13780 16244
rect 15016 16192 15068 16244
rect 16396 16192 16448 16244
rect 18512 16192 18564 16244
rect 8668 16124 8720 16176
rect 7656 15852 7708 15904
rect 8208 15852 8260 15904
rect 10600 16056 10652 16108
rect 13728 16056 13780 16108
rect 19064 16124 19116 16176
rect 20628 16167 20680 16176
rect 20628 16133 20637 16167
rect 20637 16133 20671 16167
rect 20671 16133 20680 16167
rect 20628 16124 20680 16133
rect 9404 15852 9456 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 13084 15852 13136 15904
rect 18512 16056 18564 16108
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 17776 15988 17828 16040
rect 19800 15988 19852 16040
rect 19892 15988 19944 16040
rect 18052 15963 18104 15972
rect 18052 15929 18061 15963
rect 18061 15929 18095 15963
rect 18095 15929 18104 15963
rect 18052 15920 18104 15929
rect 21272 15963 21324 15972
rect 21272 15929 21281 15963
rect 21281 15929 21315 15963
rect 21315 15929 21324 15963
rect 21272 15920 21324 15929
rect 16120 15852 16172 15904
rect 16304 15852 16356 15904
rect 19524 15852 19576 15904
rect 19892 15852 19944 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 8024 15648 8076 15700
rect 2320 15623 2372 15632
rect 2320 15589 2329 15623
rect 2329 15589 2363 15623
rect 2363 15589 2372 15623
rect 2320 15580 2372 15589
rect 10232 15648 10284 15700
rect 13452 15648 13504 15700
rect 11704 15580 11756 15632
rect 16304 15648 16356 15700
rect 16948 15691 17000 15700
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 17224 15648 17276 15700
rect 20352 15648 20404 15700
rect 5080 15555 5132 15564
rect 5080 15521 5089 15555
rect 5089 15521 5123 15555
rect 5123 15521 5132 15555
rect 5080 15512 5132 15521
rect 7196 15512 7248 15564
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 8484 15512 8536 15564
rect 8760 15512 8812 15564
rect 10600 15512 10652 15564
rect 18512 15555 18564 15564
rect 4620 15444 4672 15496
rect 6552 15487 6604 15496
rect 3056 15376 3108 15428
rect 2872 15308 2924 15360
rect 3240 15308 3292 15360
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 9220 15487 9272 15496
rect 6644 15376 6696 15428
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 8208 15308 8260 15360
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 10784 15444 10836 15496
rect 9312 15376 9364 15428
rect 10968 15376 11020 15428
rect 13268 15444 13320 15496
rect 14464 15444 14516 15496
rect 18512 15521 18521 15555
rect 18521 15521 18555 15555
rect 18555 15521 18564 15555
rect 18512 15512 18564 15521
rect 16948 15444 17000 15496
rect 20720 15487 20772 15496
rect 17040 15376 17092 15428
rect 15384 15308 15436 15360
rect 15844 15308 15896 15360
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 18328 15308 18380 15360
rect 19524 15308 19576 15360
rect 20444 15308 20496 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 3332 15104 3384 15156
rect 4068 15104 4120 15156
rect 5448 15104 5500 15156
rect 2412 15036 2464 15088
rect 8484 15036 8536 15088
rect 8760 15104 8812 15156
rect 13268 15104 13320 15156
rect 14832 15147 14884 15156
rect 14832 15113 14841 15147
rect 14841 15113 14875 15147
rect 14875 15113 14884 15147
rect 14832 15104 14884 15113
rect 15936 15147 15988 15156
rect 15476 15036 15528 15088
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 6000 14968 6052 15020
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5264 14900 5316 14909
rect 5540 14900 5592 14952
rect 6552 14900 6604 14952
rect 4712 14832 4764 14884
rect 9220 14968 9272 15020
rect 9772 14968 9824 15020
rect 10416 14968 10468 15020
rect 13544 14968 13596 15020
rect 15936 15113 15945 15147
rect 15945 15113 15979 15147
rect 15979 15113 15988 15147
rect 15936 15104 15988 15113
rect 16948 15104 17000 15156
rect 18696 15036 18748 15088
rect 17224 14968 17276 15020
rect 7840 14900 7892 14952
rect 2780 14764 2832 14816
rect 3332 14807 3384 14816
rect 3332 14773 3341 14807
rect 3341 14773 3375 14807
rect 3375 14773 3384 14807
rect 3332 14764 3384 14773
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 4436 14764 4488 14816
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7196 14764 7248 14816
rect 15476 14900 15528 14952
rect 16212 14900 16264 14952
rect 10876 14832 10928 14884
rect 13452 14832 13504 14884
rect 10324 14764 10376 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 11244 14764 11296 14816
rect 11704 14764 11756 14816
rect 13268 14764 13320 14816
rect 15752 14764 15804 14816
rect 16948 14764 17000 14816
rect 17316 14764 17368 14816
rect 18328 14764 18380 14816
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 20812 14764 20864 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 4988 14560 5040 14612
rect 5172 14560 5224 14612
rect 9772 14560 9824 14612
rect 10876 14560 10928 14612
rect 10968 14560 11020 14612
rect 13728 14560 13780 14612
rect 3792 14492 3844 14544
rect 3976 14492 4028 14544
rect 3976 14356 4028 14408
rect 4252 14424 4304 14476
rect 5080 14424 5132 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 9128 14492 9180 14544
rect 11244 14492 11296 14544
rect 11980 14492 12032 14544
rect 13452 14492 13504 14544
rect 15476 14560 15528 14612
rect 15660 14560 15712 14612
rect 16396 14560 16448 14612
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 18788 14560 18840 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 9220 14424 9272 14476
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 8392 14356 8444 14408
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 2780 14220 2832 14272
rect 5172 14288 5224 14340
rect 5632 14288 5684 14340
rect 4068 14220 4120 14272
rect 5724 14220 5776 14272
rect 6828 14220 6880 14272
rect 8392 14220 8444 14272
rect 8944 14356 8996 14408
rect 10140 14356 10192 14408
rect 10508 14399 10560 14408
rect 10508 14365 10542 14399
rect 10542 14365 10560 14399
rect 10508 14356 10560 14365
rect 9312 14288 9364 14340
rect 9496 14288 9548 14340
rect 8760 14220 8812 14272
rect 9956 14220 10008 14272
rect 10048 14220 10100 14272
rect 13544 14356 13596 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 16028 14399 16080 14408
rect 16028 14365 16062 14399
rect 16062 14365 16080 14399
rect 16028 14356 16080 14365
rect 15844 14288 15896 14340
rect 11796 14220 11848 14272
rect 12900 14220 12952 14272
rect 13544 14220 13596 14272
rect 14464 14220 14516 14272
rect 18328 14220 18380 14272
rect 19340 14356 19392 14408
rect 19524 14356 19576 14408
rect 20628 14399 20680 14408
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 20720 14356 20772 14408
rect 21272 14356 21324 14408
rect 19984 14288 20036 14340
rect 20352 14331 20404 14340
rect 20352 14297 20370 14331
rect 20370 14297 20404 14331
rect 20352 14288 20404 14297
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 5264 14016 5316 14068
rect 4068 13948 4120 14000
rect 4344 13991 4396 14000
rect 4344 13957 4353 13991
rect 4353 13957 4387 13991
rect 4387 13957 4396 13991
rect 4344 13948 4396 13957
rect 5816 13948 5868 14000
rect 8760 13948 8812 14000
rect 12808 14016 12860 14068
rect 15292 14016 15344 14068
rect 16028 14016 16080 14068
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 19708 14016 19760 14068
rect 2596 13880 2648 13932
rect 3792 13880 3844 13932
rect 8944 13880 8996 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9496 13923 9548 13932
rect 9496 13889 9530 13923
rect 9530 13889 9548 13923
rect 9496 13880 9548 13889
rect 10048 13880 10100 13932
rect 5080 13812 5132 13864
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 11796 13880 11848 13932
rect 20628 13948 20680 14000
rect 17224 13880 17276 13932
rect 17592 13923 17644 13932
rect 4068 13744 4120 13796
rect 7472 13744 7524 13796
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 12900 13855 12952 13864
rect 11704 13812 11756 13821
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 5724 13676 5776 13728
rect 10140 13676 10192 13728
rect 14464 13676 14516 13728
rect 15752 13812 15804 13864
rect 16028 13812 16080 13864
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 18328 13880 18380 13932
rect 19708 13880 19760 13932
rect 20996 13923 21048 13932
rect 20996 13889 21014 13923
rect 21014 13889 21048 13923
rect 20996 13880 21048 13889
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 1860 13472 1912 13524
rect 3424 13472 3476 13524
rect 6000 13472 6052 13524
rect 8116 13472 8168 13524
rect 6552 13404 6604 13456
rect 10508 13472 10560 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 17040 13472 17092 13524
rect 17592 13472 17644 13524
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 14556 13404 14608 13456
rect 7012 13336 7064 13345
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6828 13268 6880 13320
rect 2044 13175 2096 13184
rect 2044 13141 2053 13175
rect 2053 13141 2087 13175
rect 2087 13141 2096 13175
rect 2044 13132 2096 13141
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 2504 13132 2556 13184
rect 5448 13200 5500 13252
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 4436 13132 4488 13184
rect 5816 13132 5868 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7748 13132 7800 13184
rect 8116 13132 8168 13184
rect 9220 13336 9272 13388
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 9220 13200 9272 13252
rect 9864 13200 9916 13252
rect 12256 13200 12308 13252
rect 16396 13200 16448 13252
rect 10048 13132 10100 13184
rect 11704 13132 11756 13184
rect 17132 13132 17184 13184
rect 17316 13132 17368 13184
rect 18144 13132 18196 13184
rect 20168 13200 20220 13252
rect 20812 13200 20864 13252
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2044 12928 2096 12980
rect 4252 12928 4304 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 6184 12928 6236 12980
rect 6736 12928 6788 12980
rect 7380 12928 7432 12980
rect 8576 12928 8628 12980
rect 9312 12928 9364 12980
rect 9956 12928 10008 12980
rect 10416 12928 10468 12980
rect 10876 12928 10928 12980
rect 11704 12928 11756 12980
rect 4344 12860 4396 12912
rect 4804 12860 4856 12912
rect 8116 12860 8168 12912
rect 10232 12860 10284 12912
rect 13912 12928 13964 12980
rect 1676 12792 1728 12844
rect 2688 12792 2740 12844
rect 4988 12792 5040 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 4620 12724 4672 12776
rect 4804 12724 4856 12776
rect 6092 12792 6144 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 6000 12724 6052 12776
rect 7748 12767 7800 12776
rect 3976 12656 4028 12708
rect 4344 12656 4396 12708
rect 5632 12656 5684 12708
rect 4252 12588 4304 12640
rect 5264 12588 5316 12640
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 10876 12792 10928 12844
rect 15660 12860 15712 12912
rect 6736 12656 6788 12708
rect 14464 12792 14516 12844
rect 15752 12792 15804 12844
rect 16028 12928 16080 12980
rect 19064 12928 19116 12980
rect 19524 12928 19576 12980
rect 20168 12928 20220 12980
rect 20260 12928 20312 12980
rect 19708 12903 19760 12912
rect 19708 12869 19717 12903
rect 19717 12869 19751 12903
rect 19751 12869 19760 12903
rect 19708 12860 19760 12869
rect 17592 12792 17644 12844
rect 19800 12792 19852 12844
rect 20260 12792 20312 12844
rect 21272 12792 21324 12844
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 8208 12588 8260 12640
rect 9312 12588 9364 12640
rect 10232 12588 10284 12640
rect 19984 12656 20036 12708
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 13912 12588 13964 12640
rect 15292 12588 15344 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 4160 12384 4212 12436
rect 5632 12384 5684 12436
rect 5908 12384 5960 12436
rect 6828 12384 6880 12436
rect 3056 12316 3108 12368
rect 11796 12384 11848 12436
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 17592 12384 17644 12436
rect 20352 12384 20404 12436
rect 20996 12384 21048 12436
rect 2688 12248 2740 12300
rect 4068 12248 4120 12300
rect 6828 12248 6880 12300
rect 8668 12316 8720 12368
rect 9128 12316 9180 12368
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 2780 12180 2832 12232
rect 5908 12180 5960 12232
rect 6184 12180 6236 12232
rect 8116 12180 8168 12232
rect 13176 12316 13228 12368
rect 15660 12316 15712 12368
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 20812 12248 20864 12300
rect 1768 12112 1820 12164
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 2044 12044 2096 12096
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 2688 12044 2740 12096
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 3516 12044 3568 12096
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4896 12087 4948 12096
rect 4344 12044 4396 12053
rect 4896 12053 4905 12087
rect 4905 12053 4939 12087
rect 4939 12053 4948 12087
rect 4896 12044 4948 12053
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 6920 12044 6972 12096
rect 7104 12044 7156 12096
rect 7564 12044 7616 12096
rect 8208 12044 8260 12096
rect 10324 12155 10376 12164
rect 10324 12121 10342 12155
rect 10342 12121 10376 12155
rect 13820 12180 13872 12232
rect 14924 12180 14976 12232
rect 15752 12180 15804 12232
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 10324 12112 10376 12121
rect 13268 12112 13320 12164
rect 15292 12112 15344 12164
rect 17592 12112 17644 12164
rect 19708 12112 19760 12164
rect 19892 12112 19944 12164
rect 16948 12044 17000 12096
rect 17224 12044 17276 12096
rect 18144 12044 18196 12096
rect 18512 12044 18564 12096
rect 19616 12087 19668 12096
rect 19616 12053 19625 12087
rect 19625 12053 19659 12087
rect 19659 12053 19668 12087
rect 19616 12044 19668 12053
rect 19984 12044 20036 12096
rect 20996 12044 21048 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 2136 11840 2188 11892
rect 3240 11840 3292 11892
rect 3516 11883 3568 11892
rect 3516 11849 3525 11883
rect 3525 11849 3559 11883
rect 3559 11849 3568 11883
rect 3516 11840 3568 11849
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 4344 11840 4396 11892
rect 6644 11840 6696 11892
rect 7104 11840 7156 11892
rect 7472 11840 7524 11892
rect 7656 11840 7708 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 1860 11772 1912 11824
rect 5724 11772 5776 11824
rect 6552 11772 6604 11824
rect 7932 11772 7984 11824
rect 8208 11772 8260 11824
rect 8668 11815 8720 11824
rect 8668 11781 8677 11815
rect 8677 11781 8711 11815
rect 8711 11781 8720 11815
rect 11704 11840 11756 11892
rect 13176 11883 13228 11892
rect 8668 11772 8720 11781
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 4988 11704 5040 11756
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 2136 11500 2188 11552
rect 2688 11500 2740 11552
rect 5264 11636 5316 11688
rect 6828 11704 6880 11756
rect 11152 11772 11204 11824
rect 11612 11772 11664 11824
rect 11888 11772 11940 11824
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 5632 11568 5684 11620
rect 6092 11636 6144 11688
rect 10140 11704 10192 11756
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 13820 11772 13872 11824
rect 14832 11772 14884 11824
rect 16304 11840 16356 11892
rect 18604 11840 18656 11892
rect 20168 11840 20220 11892
rect 20628 11840 20680 11892
rect 13452 11704 13504 11756
rect 18052 11704 18104 11756
rect 19064 11772 19116 11824
rect 20260 11772 20312 11824
rect 20444 11747 20496 11756
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 17868 11636 17920 11688
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 20720 11636 20772 11688
rect 4620 11500 4672 11552
rect 6092 11500 6144 11552
rect 6552 11500 6604 11552
rect 8116 11500 8168 11552
rect 8484 11500 8536 11552
rect 11612 11568 11664 11620
rect 19800 11568 19852 11620
rect 20536 11568 20588 11620
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 20720 11500 20772 11552
rect 20996 11500 21048 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2872 11296 2924 11348
rect 5632 11296 5684 11348
rect 9956 11296 10008 11348
rect 1492 11160 1544 11212
rect 3056 11228 3108 11280
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 3148 11160 3200 11212
rect 5264 11160 5316 11212
rect 6828 11160 6880 11212
rect 6920 11160 6972 11212
rect 9404 11228 9456 11280
rect 10876 11296 10928 11348
rect 17224 11296 17276 11348
rect 19616 11296 19668 11348
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 10784 11228 10836 11280
rect 1400 11092 1452 11144
rect 3516 11092 3568 11144
rect 7932 11092 7984 11144
rect 8668 11092 8720 11144
rect 2412 11024 2464 11076
rect 4344 11067 4396 11076
rect 4344 11033 4353 11067
rect 4353 11033 4387 11067
rect 4387 11033 4396 11067
rect 4344 11024 4396 11033
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 2780 10999 2832 11008
rect 2780 10965 2789 10999
rect 2789 10965 2823 10999
rect 2823 10965 2832 10999
rect 5448 11024 5500 11076
rect 7288 11024 7340 11076
rect 8484 11024 8536 11076
rect 12072 11160 12124 11212
rect 13452 11160 13504 11212
rect 9496 11092 9548 11144
rect 13820 11092 13872 11144
rect 9680 11024 9732 11076
rect 10692 11024 10744 11076
rect 16672 11092 16724 11144
rect 17868 11092 17920 11144
rect 20628 11092 20680 11144
rect 17408 11024 17460 11076
rect 2780 10956 2832 10965
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 19892 11024 19944 11076
rect 20812 11024 20864 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2872 10752 2924 10804
rect 3424 10752 3476 10804
rect 2780 10684 2832 10736
rect 3976 10752 4028 10804
rect 6000 10752 6052 10804
rect 6644 10752 6696 10804
rect 2412 10616 2464 10668
rect 5356 10684 5408 10736
rect 9312 10752 9364 10804
rect 2136 10548 2188 10600
rect 3056 10548 3108 10600
rect 5448 10616 5500 10668
rect 5080 10548 5132 10600
rect 8576 10616 8628 10668
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 7288 10548 7340 10600
rect 7748 10548 7800 10600
rect 9956 10684 10008 10736
rect 12164 10684 12216 10736
rect 2964 10480 3016 10532
rect 6552 10480 6604 10532
rect 8668 10480 8720 10532
rect 10692 10616 10744 10668
rect 12440 10616 12492 10668
rect 14924 10616 14976 10668
rect 15200 10752 15252 10804
rect 16028 10752 16080 10804
rect 17684 10752 17736 10804
rect 19616 10752 19668 10804
rect 20628 10752 20680 10804
rect 18052 10684 18104 10736
rect 19800 10727 19852 10736
rect 19800 10693 19834 10727
rect 19834 10693 19852 10727
rect 19800 10684 19852 10693
rect 17132 10616 17184 10668
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 13820 10548 13872 10600
rect 19524 10591 19576 10600
rect 19524 10557 19533 10591
rect 19533 10557 19567 10591
rect 19567 10557 19576 10591
rect 19524 10548 19576 10557
rect 20812 10480 20864 10532
rect 4804 10412 4856 10464
rect 5540 10412 5592 10464
rect 6092 10412 6144 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 9680 10412 9732 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2872 10208 2924 10260
rect 6552 10208 6604 10260
rect 7104 10208 7156 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 2872 10115 2924 10124
rect 2872 10081 2881 10115
rect 2881 10081 2915 10115
rect 2915 10081 2924 10115
rect 2872 10072 2924 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5448 10072 5500 10124
rect 7656 10072 7708 10124
rect 9404 10208 9456 10260
rect 9956 10208 10008 10260
rect 10324 10208 10376 10260
rect 14464 10208 14516 10260
rect 17040 10208 17092 10260
rect 14556 10140 14608 10192
rect 17960 10208 18012 10260
rect 20076 10208 20128 10260
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4712 10004 4764 10056
rect 7748 10004 7800 10056
rect 9680 10004 9732 10056
rect 16396 10072 16448 10124
rect 20076 10072 20128 10124
rect 20352 10072 20404 10124
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 2964 9868 3016 9920
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4804 9868 4856 9920
rect 8024 9936 8076 9988
rect 9312 9979 9364 9988
rect 8576 9868 8628 9920
rect 9312 9945 9346 9979
rect 9346 9945 9364 9979
rect 9312 9936 9364 9945
rect 11152 9936 11204 9988
rect 13820 10004 13872 10056
rect 15752 10004 15804 10056
rect 17868 10004 17920 10056
rect 19524 10004 19576 10056
rect 16948 9979 17000 9988
rect 16948 9945 16957 9979
rect 16957 9945 16991 9979
rect 16991 9945 17000 9979
rect 16948 9936 17000 9945
rect 10784 9868 10836 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 17132 9868 17184 9920
rect 20076 9911 20128 9920
rect 20076 9877 20085 9911
rect 20085 9877 20119 9911
rect 20119 9877 20128 9911
rect 20076 9868 20128 9877
rect 20628 9868 20680 9920
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 2872 9664 2924 9716
rect 4160 9664 4212 9716
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 14464 9664 14516 9716
rect 20904 9664 20956 9716
rect 1400 9639 1452 9648
rect 1400 9605 1409 9639
rect 1409 9605 1443 9639
rect 1443 9605 1452 9639
rect 1400 9596 1452 9605
rect 3148 9596 3200 9648
rect 6000 9596 6052 9648
rect 6368 9596 6420 9648
rect 8208 9596 8260 9648
rect 9128 9596 9180 9648
rect 9404 9596 9456 9648
rect 10048 9639 10100 9648
rect 10048 9605 10082 9639
rect 10082 9605 10100 9639
rect 10048 9596 10100 9605
rect 10416 9596 10468 9648
rect 10876 9596 10928 9648
rect 17040 9596 17092 9648
rect 19616 9596 19668 9648
rect 20536 9596 20588 9648
rect 2872 9460 2924 9512
rect 3056 9460 3108 9512
rect 5540 9571 5592 9580
rect 3608 9435 3660 9444
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 3884 9392 3936 9444
rect 2964 9324 3016 9376
rect 3240 9324 3292 9376
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 5724 9528 5776 9580
rect 6092 9528 6144 9580
rect 6276 9528 6328 9580
rect 6552 9528 6604 9580
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 4528 9392 4580 9444
rect 6736 9460 6788 9512
rect 12440 9528 12492 9580
rect 9680 9460 9732 9512
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 6092 9324 6144 9376
rect 6368 9324 6420 9376
rect 6644 9324 6696 9376
rect 8484 9392 8536 9444
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 11612 9435 11664 9444
rect 11612 9401 11621 9435
rect 11621 9401 11655 9435
rect 11655 9401 11664 9435
rect 11612 9392 11664 9401
rect 9956 9324 10008 9376
rect 10508 9324 10560 9376
rect 15568 9528 15620 9580
rect 16396 9528 16448 9580
rect 17960 9528 18012 9580
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 20352 9528 20404 9580
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 21272 9528 21324 9580
rect 19708 9460 19760 9469
rect 16212 9324 16264 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1860 9120 1912 9172
rect 3240 9120 3292 9172
rect 4068 9120 4120 9172
rect 6000 9120 6052 9172
rect 7288 9120 7340 9172
rect 9772 9120 9824 9172
rect 10048 9120 10100 9172
rect 1400 9052 1452 9104
rect 3332 8984 3384 9036
rect 3884 9027 3936 9036
rect 3884 8993 3893 9027
rect 3893 8993 3927 9027
rect 3927 8993 3936 9027
rect 3884 8984 3936 8993
rect 9312 9052 9364 9104
rect 3056 8916 3108 8968
rect 4436 8916 4488 8968
rect 5632 8984 5684 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 8024 8984 8076 9036
rect 9036 8984 9088 9036
rect 10416 8984 10468 9036
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 13268 9120 13320 9172
rect 13728 9120 13780 9172
rect 14280 9120 14332 9172
rect 17684 9120 17736 9172
rect 19616 9120 19668 9172
rect 17868 9052 17920 9104
rect 19800 9052 19852 9104
rect 20168 9052 20220 9104
rect 20536 9052 20588 9104
rect 5724 8916 5776 8968
rect 5908 8916 5960 8968
rect 8668 8916 8720 8968
rect 9956 8916 10008 8968
rect 10232 8916 10284 8968
rect 10968 8916 11020 8968
rect 11612 8916 11664 8968
rect 2964 8848 3016 8900
rect 1400 8780 1452 8832
rect 3240 8780 3292 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 5724 8780 5776 8832
rect 5908 8780 5960 8832
rect 6920 8848 6972 8900
rect 8484 8848 8536 8900
rect 9772 8848 9824 8900
rect 10416 8848 10468 8900
rect 17040 8984 17092 9036
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 6460 8780 6512 8832
rect 6644 8780 6696 8832
rect 7104 8780 7156 8832
rect 7656 8780 7708 8832
rect 11796 8780 11848 8832
rect 13728 8916 13780 8968
rect 15384 8916 15436 8968
rect 15844 8916 15896 8968
rect 16028 8959 16080 8968
rect 16028 8925 16062 8959
rect 16062 8925 16080 8959
rect 16028 8916 16080 8925
rect 13268 8848 13320 8900
rect 15660 8848 15712 8900
rect 17960 8848 18012 8900
rect 14924 8780 14976 8832
rect 17040 8780 17092 8832
rect 17224 8780 17276 8832
rect 17408 8780 17460 8832
rect 19616 8916 19668 8968
rect 20260 8916 20312 8968
rect 18788 8848 18840 8900
rect 18880 8780 18932 8832
rect 20536 8780 20588 8832
rect 20812 8780 20864 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1768 8576 1820 8628
rect 1952 8576 2004 8628
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 4896 8576 4948 8628
rect 5540 8619 5592 8628
rect 2872 8508 2924 8560
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 7840 8576 7892 8628
rect 8208 8576 8260 8628
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2872 8372 2924 8424
rect 15108 8576 15160 8628
rect 8668 8508 8720 8560
rect 9496 8508 9548 8560
rect 14924 8508 14976 8560
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4712 8440 4764 8492
rect 6920 8440 6972 8492
rect 8484 8440 8536 8492
rect 14464 8440 14516 8492
rect 17132 8576 17184 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18972 8576 19024 8628
rect 19064 8508 19116 8560
rect 5080 8372 5132 8424
rect 5264 8372 5316 8424
rect 2136 8304 2188 8356
rect 7288 8372 7340 8424
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 9220 8372 9272 8424
rect 13268 8372 13320 8424
rect 13360 8372 13412 8424
rect 14280 8372 14332 8424
rect 15844 8372 15896 8424
rect 19708 8440 19760 8492
rect 9036 8304 9088 8356
rect 11796 8304 11848 8356
rect 9220 8236 9272 8288
rect 10232 8236 10284 8288
rect 10600 8236 10652 8288
rect 12164 8236 12216 8288
rect 13636 8279 13688 8288
rect 13636 8245 13645 8279
rect 13645 8245 13679 8279
rect 13679 8245 13688 8279
rect 13636 8236 13688 8245
rect 15108 8236 15160 8288
rect 18236 8304 18288 8356
rect 19800 8347 19852 8356
rect 19800 8313 19809 8347
rect 19809 8313 19843 8347
rect 19843 8313 19852 8347
rect 19800 8304 19852 8313
rect 15844 8279 15896 8288
rect 15844 8245 15853 8279
rect 15853 8245 15887 8279
rect 15887 8245 15896 8279
rect 15844 8236 15896 8245
rect 16396 8236 16448 8288
rect 17408 8236 17460 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 2412 8032 2464 8084
rect 3976 8032 4028 8084
rect 5080 8032 5132 8084
rect 6000 8032 6052 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 9588 8032 9640 8084
rect 12164 8032 12216 8084
rect 17960 8075 18012 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 3148 7964 3200 8016
rect 4068 7964 4120 8016
rect 2412 7828 2464 7880
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 1584 7760 1636 7812
rect 3976 7896 4028 7948
rect 6552 7964 6604 8016
rect 7012 7964 7064 8016
rect 5724 7939 5776 7948
rect 3240 7828 3292 7880
rect 3516 7828 3568 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 15292 7896 15344 7948
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 18328 8032 18380 8084
rect 20444 8032 20496 8084
rect 20996 8075 21048 8084
rect 20996 8041 21005 8075
rect 21005 8041 21039 8075
rect 21039 8041 21048 8075
rect 20996 8032 21048 8041
rect 19064 7964 19116 8016
rect 18052 7896 18104 7948
rect 20260 7964 20312 8016
rect 20536 7939 20588 7948
rect 9220 7828 9272 7880
rect 9312 7828 9364 7880
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3424 7760 3476 7812
rect 5264 7692 5316 7744
rect 5724 7692 5776 7744
rect 6000 7692 6052 7744
rect 6552 7692 6604 7744
rect 8668 7760 8720 7812
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 8484 7692 8536 7744
rect 10232 7828 10284 7880
rect 11152 7828 11204 7880
rect 11704 7692 11756 7744
rect 15660 7828 15712 7880
rect 16120 7871 16172 7880
rect 16120 7837 16143 7871
rect 16143 7837 16172 7871
rect 16120 7828 16172 7837
rect 17408 7828 17460 7880
rect 19984 7828 20036 7880
rect 20260 7828 20312 7880
rect 20536 7905 20545 7939
rect 20545 7905 20579 7939
rect 20579 7905 20588 7939
rect 20536 7896 20588 7905
rect 14464 7760 14516 7812
rect 17316 7692 17368 7744
rect 19984 7692 20036 7744
rect 20444 7692 20496 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 4068 7488 4120 7540
rect 4896 7488 4948 7540
rect 6000 7531 6052 7540
rect 6000 7497 6009 7531
rect 6009 7497 6043 7531
rect 6043 7497 6052 7531
rect 6000 7488 6052 7497
rect 8208 7488 8260 7540
rect 10784 7488 10836 7540
rect 17592 7488 17644 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 3240 7420 3292 7472
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 7288 7420 7340 7472
rect 10600 7420 10652 7472
rect 10692 7420 10744 7472
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2688 7284 2740 7336
rect 2780 7284 2832 7336
rect 3976 7284 4028 7336
rect 4068 7284 4120 7336
rect 7196 7352 7248 7404
rect 9220 7352 9272 7404
rect 13452 7352 13504 7404
rect 18972 7420 19024 7472
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 5632 7216 5684 7268
rect 9772 7216 9824 7268
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 7564 7148 7616 7200
rect 7840 7148 7892 7200
rect 9128 7148 9180 7200
rect 10048 7148 10100 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11152 7148 11204 7200
rect 15292 7259 15344 7268
rect 13636 7148 13688 7200
rect 15292 7225 15301 7259
rect 15301 7225 15335 7259
rect 15335 7225 15344 7259
rect 15292 7216 15344 7225
rect 17960 7352 18012 7404
rect 18328 7395 18380 7404
rect 18328 7361 18337 7395
rect 18337 7361 18371 7395
rect 18371 7361 18380 7395
rect 18328 7352 18380 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 21180 7352 21232 7404
rect 19064 7284 19116 7336
rect 20076 7284 20128 7336
rect 16304 7216 16356 7268
rect 18420 7216 18472 7268
rect 20352 7216 20404 7268
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15568 7148 15620 7200
rect 16396 7148 16448 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2228 6944 2280 6996
rect 7012 6944 7064 6996
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 3424 6876 3476 6928
rect 4068 6876 4120 6928
rect 5080 6808 5132 6860
rect 6000 6808 6052 6860
rect 7564 6876 7616 6928
rect 18420 6944 18472 6996
rect 19064 6944 19116 6996
rect 6828 6808 6880 6860
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 17960 6876 18012 6928
rect 18328 6876 18380 6928
rect 18604 6876 18656 6928
rect 8024 6808 8076 6817
rect 3148 6740 3200 6792
rect 3424 6740 3476 6792
rect 4896 6740 4948 6792
rect 5356 6740 5408 6792
rect 6920 6740 6972 6792
rect 7104 6740 7156 6792
rect 7472 6740 7524 6792
rect 9772 6740 9824 6792
rect 20076 6808 20128 6860
rect 20352 6808 20404 6860
rect 11060 6740 11112 6792
rect 1768 6672 1820 6724
rect 5816 6672 5868 6724
rect 3056 6604 3108 6656
rect 3240 6604 3292 6656
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 7012 6604 7064 6656
rect 8484 6672 8536 6724
rect 10508 6672 10560 6724
rect 11980 6740 12032 6792
rect 13636 6740 13688 6792
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 18880 6740 18932 6792
rect 20168 6740 20220 6792
rect 11244 6672 11296 6724
rect 16028 6672 16080 6724
rect 18512 6672 18564 6724
rect 18788 6715 18840 6724
rect 18788 6681 18797 6715
rect 18797 6681 18831 6715
rect 18831 6681 18840 6715
rect 18788 6672 18840 6681
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 9128 6604 9180 6656
rect 9404 6604 9456 6656
rect 11060 6604 11112 6656
rect 11704 6604 11756 6656
rect 15752 6604 15804 6656
rect 17132 6604 17184 6656
rect 18236 6604 18288 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 18604 6604 18656 6656
rect 19524 6604 19576 6656
rect 19616 6604 19668 6656
rect 20812 6672 20864 6724
rect 21364 6672 21416 6724
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 20904 6604 20956 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 1952 6400 2004 6452
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 2964 6400 3016 6452
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5264 6400 5316 6452
rect 9588 6400 9640 6452
rect 13452 6443 13504 6452
rect 13452 6409 13461 6443
rect 13461 6409 13495 6443
rect 13495 6409 13504 6443
rect 13452 6400 13504 6409
rect 15476 6400 15528 6452
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 17960 6400 18012 6452
rect 7012 6332 7064 6384
rect 7748 6332 7800 6384
rect 8852 6332 8904 6384
rect 15936 6375 15988 6384
rect 15936 6341 15945 6375
rect 15945 6341 15979 6375
rect 15979 6341 15988 6375
rect 15936 6332 15988 6341
rect 1400 6264 1452 6316
rect 2688 6264 2740 6316
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 6920 6307 6972 6316
rect 1768 6196 1820 6248
rect 1584 6128 1636 6180
rect 2320 6196 2372 6248
rect 3976 6196 4028 6248
rect 6000 6196 6052 6248
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 8576 6307 8628 6316
rect 7564 6264 7616 6273
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 9404 6264 9456 6316
rect 12164 6264 12216 6316
rect 16120 6264 16172 6316
rect 17040 6307 17092 6316
rect 7104 6196 7156 6248
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 2964 6060 3016 6112
rect 4528 6060 4580 6112
rect 5080 6060 5132 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 5632 6060 5684 6112
rect 6828 6060 6880 6112
rect 8852 6196 8904 6248
rect 8944 6171 8996 6180
rect 8944 6137 8953 6171
rect 8953 6137 8987 6171
rect 8987 6137 8996 6171
rect 8944 6128 8996 6137
rect 9680 6128 9732 6180
rect 9404 6060 9456 6112
rect 11704 6196 11756 6248
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 16396 6196 16448 6248
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 19708 6332 19760 6384
rect 18236 6264 18288 6316
rect 19064 6264 19116 6316
rect 17776 6128 17828 6180
rect 13452 6060 13504 6112
rect 13636 6060 13688 6112
rect 18236 6128 18288 6180
rect 18696 6196 18748 6248
rect 19616 6264 19668 6316
rect 20076 6307 20128 6316
rect 20076 6273 20094 6307
rect 20094 6273 20128 6307
rect 20076 6264 20128 6273
rect 20352 6307 20404 6316
rect 20352 6273 20361 6307
rect 20361 6273 20395 6307
rect 20395 6273 20404 6307
rect 20996 6307 21048 6316
rect 20352 6264 20404 6273
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 18972 6128 19024 6180
rect 21364 6264 21416 6316
rect 18144 6060 18196 6112
rect 20904 6060 20956 6112
rect 21088 6060 21140 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 4068 5856 4120 5908
rect 4620 5856 4672 5908
rect 5356 5856 5408 5908
rect 5540 5856 5592 5908
rect 7380 5856 7432 5908
rect 4528 5788 4580 5840
rect 1676 5720 1728 5772
rect 3148 5763 3200 5772
rect 3148 5729 3157 5763
rect 3157 5729 3191 5763
rect 3191 5729 3200 5763
rect 3148 5720 3200 5729
rect 3976 5720 4028 5772
rect 6000 5788 6052 5840
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 7472 5720 7524 5772
rect 9312 5788 9364 5840
rect 11980 5856 12032 5908
rect 18604 5856 18656 5908
rect 5448 5652 5500 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 7564 5584 7616 5636
rect 1768 5516 1820 5568
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 6736 5516 6788 5568
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8668 5584 8720 5636
rect 9956 5584 10008 5636
rect 10048 5584 10100 5636
rect 9312 5516 9364 5568
rect 10232 5516 10284 5568
rect 11244 5516 11296 5568
rect 13452 5720 13504 5772
rect 20352 5856 20404 5908
rect 20628 5856 20680 5908
rect 15568 5695 15620 5704
rect 12440 5584 12492 5636
rect 14464 5584 14516 5636
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 18236 5652 18288 5704
rect 21180 5788 21232 5840
rect 17224 5627 17276 5636
rect 17224 5593 17242 5627
rect 17242 5593 17276 5627
rect 17224 5584 17276 5593
rect 17684 5584 17736 5636
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 13820 5516 13872 5568
rect 15752 5516 15804 5568
rect 18052 5516 18104 5568
rect 19156 5516 19208 5568
rect 19708 5516 19760 5568
rect 20168 5516 20220 5568
rect 20536 5516 20588 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2596 5355 2648 5364
rect 2596 5321 2605 5355
rect 2605 5321 2639 5355
rect 2639 5321 2648 5355
rect 2596 5312 2648 5321
rect 3148 5312 3200 5364
rect 4160 5312 4212 5364
rect 5264 5312 5316 5364
rect 6828 5312 6880 5364
rect 9220 5312 9272 5364
rect 13728 5312 13780 5364
rect 4620 5244 4672 5296
rect 2320 5108 2372 5160
rect 3148 5040 3200 5092
rect 1768 4972 1820 5024
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 8392 5176 8444 5228
rect 11704 5244 11756 5296
rect 10140 5176 10192 5228
rect 13728 5176 13780 5228
rect 15292 5312 15344 5364
rect 15568 5312 15620 5364
rect 16856 5312 16908 5364
rect 17500 5312 17552 5364
rect 15384 5287 15436 5296
rect 15384 5253 15393 5287
rect 15393 5253 15427 5287
rect 15427 5253 15436 5287
rect 15384 5244 15436 5253
rect 20720 5244 20772 5296
rect 20904 5287 20956 5296
rect 20904 5253 20913 5287
rect 20913 5253 20947 5287
rect 20947 5253 20956 5287
rect 20904 5244 20956 5253
rect 4620 5108 4672 5160
rect 6000 5108 6052 5160
rect 7656 5108 7708 5160
rect 16580 5176 16632 5228
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 18972 5176 19024 5228
rect 20536 5176 20588 5228
rect 3976 4972 4028 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 4896 4972 4948 5024
rect 11244 5040 11296 5092
rect 12440 5083 12492 5092
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 11704 4972 11756 5024
rect 16304 5108 16356 5160
rect 18236 5108 18288 5160
rect 15568 5040 15620 5092
rect 18144 5083 18196 5092
rect 18144 5049 18153 5083
rect 18153 5049 18187 5083
rect 18187 5049 18196 5083
rect 18144 5040 18196 5049
rect 18604 5040 18656 5092
rect 19156 5108 19208 5160
rect 19064 5040 19116 5092
rect 20812 5108 20864 5160
rect 20536 5083 20588 5092
rect 20536 5049 20545 5083
rect 20545 5049 20579 5083
rect 20579 5049 20588 5083
rect 20536 5040 20588 5049
rect 20904 4972 20956 5024
rect 21088 4972 21140 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 1676 4768 1728 4820
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 2504 4768 2556 4820
rect 7104 4768 7156 4820
rect 4712 4700 4764 4752
rect 4068 4632 4120 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 5172 4632 5224 4684
rect 1768 4564 1820 4616
rect 2412 4564 2464 4616
rect 3148 4564 3200 4616
rect 4436 4564 4488 4616
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 9772 4700 9824 4752
rect 10416 4700 10468 4752
rect 12164 4768 12216 4820
rect 16120 4768 16172 4820
rect 12624 4700 12676 4752
rect 6552 4564 6604 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 10692 4632 10744 4684
rect 13728 4632 13780 4684
rect 17316 4768 17368 4820
rect 20168 4768 20220 4820
rect 20904 4811 20956 4820
rect 20904 4777 20913 4811
rect 20913 4777 20947 4811
rect 20947 4777 20956 4811
rect 20904 4768 20956 4777
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 3976 4428 4028 4480
rect 5172 4428 5224 4480
rect 7196 4496 7248 4548
rect 11152 4496 11204 4548
rect 12164 4496 12216 4548
rect 7840 4428 7892 4480
rect 10048 4428 10100 4480
rect 15200 4471 15252 4480
rect 15200 4437 15209 4471
rect 15209 4437 15243 4471
rect 15243 4437 15252 4471
rect 15200 4428 15252 4437
rect 19800 4564 19852 4616
rect 19892 4496 19944 4548
rect 20260 4428 20312 4480
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 21364 4428 21416 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 2964 4224 3016 4276
rect 7932 4267 7984 4276
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 9128 4224 9180 4276
rect 10600 4224 10652 4276
rect 2228 4156 2280 4208
rect 4252 4156 4304 4208
rect 4620 4156 4672 4208
rect 10876 4199 10928 4208
rect 10876 4165 10894 4199
rect 10894 4165 10928 4199
rect 10876 4156 10928 4165
rect 15292 4224 15344 4276
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 2596 4088 2648 4140
rect 5908 4088 5960 4140
rect 6552 4088 6604 4140
rect 8484 4088 8536 4140
rect 8576 4088 8628 4140
rect 8944 4088 8996 4140
rect 2688 4020 2740 4072
rect 5816 4020 5868 4072
rect 7012 4020 7064 4072
rect 7288 4020 7340 4072
rect 6000 3952 6052 4004
rect 9588 4020 9640 4072
rect 11336 4088 11388 4140
rect 11704 4088 11756 4140
rect 12164 4156 12216 4208
rect 18144 4224 18196 4276
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 15292 4131 15344 4140
rect 13452 4088 13504 4097
rect 15292 4097 15310 4131
rect 15310 4097 15344 4131
rect 15292 4088 15344 4097
rect 20352 4156 20404 4208
rect 17316 4088 17368 4140
rect 19708 4088 19760 4140
rect 20628 4088 20680 4140
rect 21272 4131 21324 4140
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 9772 3995 9824 4004
rect 9772 3961 9781 3995
rect 9781 3961 9815 3995
rect 9815 3961 9824 3995
rect 9772 3952 9824 3961
rect 11152 3952 11204 4004
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 4344 3884 4396 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 7288 3884 7340 3936
rect 8484 3884 8536 3936
rect 9404 3884 9456 3936
rect 9864 3884 9916 3936
rect 11336 3884 11388 3936
rect 12072 3884 12124 3936
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14464 3884 14516 3936
rect 15292 3884 15344 3936
rect 16212 3952 16264 4004
rect 16396 3952 16448 4004
rect 17684 4063 17736 4072
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 18880 4020 18932 4072
rect 18696 3952 18748 4004
rect 18788 3952 18840 4004
rect 17960 3884 18012 3936
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2504 3680 2556 3732
rect 2688 3680 2740 3732
rect 3976 3680 4028 3732
rect 5264 3680 5316 3732
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 8852 3680 8904 3732
rect 10600 3723 10652 3732
rect 2320 3612 2372 3664
rect 5724 3612 5776 3664
rect 6736 3655 6788 3664
rect 6736 3621 6745 3655
rect 6745 3621 6779 3655
rect 6779 3621 6788 3655
rect 6736 3612 6788 3621
rect 9312 3612 9364 3664
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 10876 3680 10928 3732
rect 12532 3680 12584 3732
rect 14372 3723 14424 3732
rect 2136 3587 2188 3596
rect 2136 3553 2145 3587
rect 2145 3553 2179 3587
rect 2179 3553 2188 3587
rect 2136 3544 2188 3553
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 5540 3544 5592 3596
rect 7288 3544 7340 3596
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 4712 3476 4764 3528
rect 7012 3519 7064 3528
rect 2596 3408 2648 3460
rect 3056 3408 3108 3460
rect 2964 3340 3016 3392
rect 4804 3408 4856 3460
rect 5540 3408 5592 3460
rect 5908 3408 5960 3460
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 8116 3476 8168 3528
rect 8852 3408 8904 3460
rect 10140 3544 10192 3596
rect 12072 3612 12124 3664
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 16580 3680 16632 3732
rect 17592 3680 17644 3732
rect 17868 3723 17920 3732
rect 17868 3689 17877 3723
rect 17877 3689 17911 3723
rect 17911 3689 17920 3723
rect 17868 3680 17920 3689
rect 15568 3612 15620 3664
rect 16672 3612 16724 3664
rect 18052 3612 18104 3664
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15108 3544 15160 3596
rect 17316 3587 17368 3596
rect 12624 3476 12676 3528
rect 11612 3408 11664 3460
rect 11796 3408 11848 3460
rect 12440 3408 12492 3460
rect 13820 3476 13872 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 18236 3612 18288 3664
rect 18420 3544 18472 3596
rect 17868 3476 17920 3528
rect 17960 3476 18012 3528
rect 18880 3544 18932 3596
rect 19064 3612 19116 3664
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 20260 3476 20312 3528
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 21180 3476 21232 3528
rect 3976 3340 4028 3392
rect 6920 3340 6972 3392
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 9036 3340 9088 3392
rect 9496 3340 9548 3392
rect 16304 3340 16356 3392
rect 21364 3340 21416 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 3976 3136 4028 3188
rect 4068 3136 4120 3188
rect 3884 3068 3936 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 4252 3136 4304 3188
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5908 3136 5960 3188
rect 4988 3068 5040 3120
rect 6920 3068 6972 3120
rect 8116 3068 8168 3120
rect 9496 3068 9548 3120
rect 13268 3179 13320 3188
rect 12900 3068 12952 3120
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 13544 3136 13596 3188
rect 16304 3136 16356 3188
rect 16948 3136 17000 3188
rect 18144 3136 18196 3188
rect 18696 3136 18748 3188
rect 18972 3136 19024 3188
rect 20628 3136 20680 3188
rect 21456 3136 21508 3188
rect 7656 3043 7708 3052
rect 5172 2932 5224 2984
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 9772 3000 9824 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11704 3000 11756 3052
rect 5632 2864 5684 2916
rect 10140 2932 10192 2984
rect 2136 2839 2188 2848
rect 2136 2805 2145 2839
rect 2145 2805 2179 2839
rect 2179 2805 2188 2839
rect 2136 2796 2188 2805
rect 2964 2796 3016 2848
rect 3332 2796 3384 2848
rect 5356 2796 5408 2848
rect 5724 2796 5776 2848
rect 12440 2932 12492 2984
rect 13176 2975 13228 2984
rect 13176 2941 13185 2975
rect 13185 2941 13219 2975
rect 13219 2941 13228 2975
rect 13176 2932 13228 2941
rect 14280 3000 14332 3052
rect 14740 3000 14792 3052
rect 15752 3068 15804 3120
rect 16028 3068 16080 3120
rect 14188 2932 14240 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 15200 2932 15252 2984
rect 18604 3068 18656 3120
rect 17960 3000 18012 3052
rect 18880 3000 18932 3052
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 20628 3000 20680 3052
rect 9680 2796 9732 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 14740 2864 14792 2916
rect 15660 2864 15712 2916
rect 16212 2864 16264 2916
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 19800 2932 19852 2984
rect 9772 2796 9824 2805
rect 14280 2796 14332 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 2780 2592 2832 2644
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 11152 2592 11204 2644
rect 12440 2592 12492 2644
rect 13176 2592 13228 2644
rect 14280 2592 14332 2644
rect 2136 2524 2188 2576
rect 13268 2524 13320 2576
rect 15200 2592 15252 2644
rect 17224 2592 17276 2644
rect 20444 2592 20496 2644
rect 1676 2456 1728 2508
rect 5264 2456 5316 2508
rect 7564 2456 7616 2508
rect 8576 2456 8628 2508
rect 12164 2456 12216 2508
rect 18420 2524 18472 2576
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 15660 2456 15712 2508
rect 21180 2499 21232 2508
rect 5540 2388 5592 2440
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 4712 2320 4764 2372
rect 5632 2320 5684 2372
rect 8668 2388 8720 2440
rect 9128 2388 9180 2440
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10140 2388 10192 2440
rect 11244 2388 11296 2440
rect 9496 2320 9548 2372
rect 14372 2388 14424 2440
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15844 2388 15896 2440
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 18328 2388 18380 2440
rect 18880 2388 18932 2440
rect 20168 2388 20220 2440
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 7840 2252 7892 2304
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 8852 2252 8904 2304
rect 10140 2252 10192 2304
rect 15016 2320 15068 2372
rect 10876 2295 10928 2304
rect 10876 2261 10885 2295
rect 10885 2261 10919 2295
rect 10919 2261 10928 2295
rect 10876 2252 10928 2261
rect 15200 2252 15252 2304
rect 16948 2320 17000 2372
rect 18604 2320 18656 2372
rect 16396 2252 16448 2304
rect 17316 2252 17368 2304
rect 17684 2252 17736 2304
rect 20260 2295 20312 2304
rect 20260 2261 20269 2295
rect 20269 2261 20303 2295
rect 20303 2261 20312 2295
rect 20260 2252 20312 2261
rect 21088 2295 21140 2304
rect 21088 2261 21097 2295
rect 21097 2261 21131 2295
rect 21131 2261 21140 2295
rect 21088 2252 21140 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 8024 2048 8076 2100
rect 12532 2048 12584 2100
rect 13268 2048 13320 2100
rect 19524 2048 19576 2100
rect 10876 1980 10928 2032
rect 15844 1980 15896 2032
rect 7840 1912 7892 1964
rect 13268 1912 13320 1964
rect 10140 1844 10192 1896
rect 15108 1844 15160 1896
rect 7288 1776 7340 1828
rect 13544 1776 13596 1828
rect 9588 1640 9640 1692
rect 10508 1640 10560 1692
rect 9312 1368 9364 1420
rect 13636 1368 13688 1420
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 3330 21312 3386 21321
rect 3330 21247 3386 21256
rect 1950 20904 2006 20913
rect 1950 20839 2006 20848
rect 1964 20602 1992 20839
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 2778 20496 2834 20505
rect 2778 20431 2834 20440
rect 2792 20058 2820 20431
rect 2870 20088 2926 20097
rect 2780 20052 2832 20058
rect 2870 20023 2926 20032
rect 2780 19994 2832 20000
rect 1952 19712 2004 19718
rect 1950 19680 1952 19689
rect 2004 19680 2006 19689
rect 1950 19615 2006 19624
rect 2884 19514 2912 20023
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 1950 19272 2006 19281
rect 1950 19207 1952 19216
rect 2004 19207 2006 19216
rect 1952 19178 2004 19184
rect 1858 18864 1914 18873
rect 1858 18799 1914 18808
rect 1768 18692 1820 18698
rect 1768 18634 1820 18640
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1490 17640 1546 17649
rect 1490 17575 1546 17584
rect 1504 17338 1532 17575
rect 1492 17332 1544 17338
rect 1492 17274 1544 17280
rect 1596 17241 1624 18022
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1582 17232 1638 17241
rect 1688 17202 1716 17478
rect 1582 17167 1638 17176
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1584 17060 1636 17066
rect 1584 17002 1636 17008
rect 1596 16574 1624 17002
rect 1688 16794 1716 17138
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1780 16574 1808 18634
rect 1872 17882 1900 18799
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18057 1992 18566
rect 2412 18080 2464 18086
rect 1950 18048 2006 18057
rect 2412 18022 2464 18028
rect 1950 17983 2006 17992
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 2424 17678 2452 18022
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16658 1992 17138
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1504 16546 1624 16574
rect 1688 16546 1808 16574
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 14793 1440 15846
rect 1398 14784 1454 14793
rect 1398 14719 1454 14728
rect 1504 12186 1532 16546
rect 1688 13002 1716 16546
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 2056 16114 2084 16458
rect 2148 16425 2176 16934
rect 2134 16416 2190 16425
rect 2134 16351 2190 16360
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2320 15632 2372 15638
rect 2318 15600 2320 15609
rect 2372 15600 2374 15609
rect 2318 15535 2374 15544
rect 2424 15094 2452 17614
rect 2516 16574 2544 19314
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 17882 2820 18391
rect 3160 18222 3188 18566
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 17202 3004 17478
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2778 16824 2834 16833
rect 2778 16759 2834 16768
rect 2516 16546 2728 16574
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 13569 1808 13670
rect 1766 13560 1822 13569
rect 1872 13530 1900 14962
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1766 13495 1822 13504
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1964 13161 1992 14214
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2044 13184 2096 13190
rect 1950 13152 2006 13161
rect 2044 13126 2096 13132
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 1950 13087 2006 13096
rect 1412 12158 1532 12186
rect 1596 12974 1716 13002
rect 2056 12986 2084 13126
rect 2044 12980 2096 12986
rect 1412 11150 1440 12158
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11218 1532 12038
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 9654 1440 11086
rect 1400 9648 1452 9654
rect 1400 9590 1452 9596
rect 1412 9110 1440 9590
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 6322 1440 8774
rect 1596 8265 1624 12974
rect 2044 12922 2096 12928
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 10810 1716 12786
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1780 12170 1808 12718
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1780 11694 1808 12106
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1780 8634 1808 10950
rect 1872 9178 1900 11766
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1582 7848 1638 7857
rect 1582 7783 1584 7792
rect 1636 7783 1638 7792
rect 1584 7754 1636 7760
rect 1596 7546 1624 7754
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 6914 1716 7890
rect 1872 7750 1900 9114
rect 1964 8634 1992 12718
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11898 2084 12038
rect 2148 11898 2176 13126
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 10606 2176 11494
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2148 9382 2176 10542
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1596 6886 1716 6914
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 3942 1440 6258
rect 1596 6186 1624 6886
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6254 1808 6666
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1584 6180 1636 6186
rect 1584 6122 1636 6128
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1688 4826 1716 5714
rect 1780 5574 1808 6190
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 5030 1808 5510
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 3777 1440 3878
rect 1398 3768 1454 3777
rect 1398 3703 1454 3712
rect 1688 2514 1716 4762
rect 1780 4622 1808 4966
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1780 3942 1808 4558
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3369 1808 3878
rect 1766 3360 1822 3369
rect 1766 3295 1822 3304
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1872 2145 1900 7686
rect 1964 6458 1992 8434
rect 2148 8362 2176 9318
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2240 8090 2268 12038
rect 2332 11801 2360 13330
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2318 11792 2374 11801
rect 2318 11727 2374 11736
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2424 11082 2452 11154
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10674 2452 11018
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2332 7546 2360 9862
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2424 7886 2452 8026
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 7002 2268 7278
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2134 5400 2190 5409
rect 2134 5335 2190 5344
rect 1950 4992 2006 5001
rect 1950 4927 2006 4936
rect 1964 3058 1992 4927
rect 2148 4826 2176 5335
rect 2332 5166 2360 6190
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2228 4208 2280 4214
rect 2228 4150 2280 4156
rect 2134 4040 2190 4049
rect 2134 3975 2190 3984
rect 2148 3602 2176 3975
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2148 2582 2176 2790
rect 2136 2576 2188 2582
rect 2136 2518 2188 2524
rect 1858 2136 1914 2145
rect 1858 2071 1914 2080
rect 2240 800 2268 4150
rect 2332 3670 2360 5102
rect 2424 4622 2452 5510
rect 2516 4826 2544 13126
rect 2608 6458 2636 13874
rect 2700 12850 2728 16546
rect 2792 16250 2820 16759
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2884 16017 2912 16934
rect 2976 16561 3004 17138
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2962 16552 3018 16561
rect 2962 16487 3018 16496
rect 2870 16008 2926 16017
rect 2870 15943 2926 15952
rect 3068 15858 3096 16934
rect 3160 15994 3188 18158
rect 3252 17746 3280 18226
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3344 17270 3372 21247
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3896 17338 3924 19790
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3332 17264 3384 17270
rect 3332 17206 3384 17212
rect 3344 16794 3372 17206
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3160 15966 3280 15994
rect 3068 15830 3188 15858
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 15026 2912 15302
rect 2962 15192 3018 15201
rect 2962 15127 3018 15136
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14385 2820 14758
rect 2778 14376 2834 14385
rect 2778 14311 2834 14320
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 12102 2728 12242
rect 2792 12238 2820 14214
rect 2780 12232 2832 12238
rect 2884 12209 2912 14962
rect 2780 12174 2832 12180
rect 2870 12200 2926 12209
rect 2870 12135 2926 12144
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 11558 2728 12038
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2884 11354 2912 11630
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10742 2820 10950
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2884 10282 2912 10746
rect 2976 10538 3004 15127
rect 3068 12481 3096 15370
rect 3054 12472 3110 12481
rect 3054 12407 3110 12416
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3068 11529 3096 12310
rect 3160 11937 3188 15830
rect 3252 15366 3280 15966
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 13410 3280 15302
rect 3344 15162 3372 16730
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3344 13977 3372 14758
rect 3330 13968 3386 13977
rect 3330 13903 3386 13912
rect 3436 13530 3464 16458
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3804 13938 3832 14486
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3252 13382 3464 13410
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3146 11928 3202 11937
rect 3252 11898 3280 12038
rect 3146 11863 3202 11872
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3054 11520 3110 11529
rect 3054 11455 3110 11464
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3068 11098 3096 11222
rect 3160 11218 3188 11698
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3068 11070 3188 11098
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2792 10266 2912 10282
rect 2792 10260 2924 10266
rect 2792 10254 2872 10260
rect 2792 8514 2820 10254
rect 2872 10202 2924 10208
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 9722 2912 10066
rect 2964 9920 3016 9926
rect 3068 9908 3096 10542
rect 3016 9880 3096 9908
rect 2964 9862 3016 9868
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 8566 2912 9454
rect 2976 9382 3004 9862
rect 3160 9738 3188 11070
rect 3068 9710 3188 9738
rect 3068 9518 3096 9710
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8906 3004 9318
rect 3068 8974 3096 9454
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2700 8486 2820 8514
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2700 7342 2728 8486
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2884 7886 2912 8366
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2976 7698 3004 8842
rect 2884 7670 3004 7698
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6322 2728 7142
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2688 5568 2740 5574
rect 2594 5536 2650 5545
rect 2688 5510 2740 5516
rect 2594 5471 2650 5480
rect 2608 5370 2636 5471
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2608 4146 2636 5306
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2516 3738 2544 4082
rect 2700 4078 2728 5510
rect 2792 4593 2820 7278
rect 2778 4584 2834 4593
rect 2778 4519 2834 4528
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2700 3534 2728 3674
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2608 800 2636 3402
rect 2792 2650 2820 4422
rect 2884 4185 2912 7670
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6458 3004 7142
rect 3068 6662 3096 8910
rect 3160 8650 3188 9590
rect 3252 9382 3280 11834
rect 3436 10810 3464 13382
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11898 3556 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3528 10554 3556 11086
rect 3344 10526 3556 10554
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9178 3280 9318
rect 3344 9217 3372 10526
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3896 10169 3924 16730
rect 3988 16182 4016 19246
rect 4080 18290 4108 20198
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4724 19514 4752 19790
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5092 18970 5120 19314
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 17338 4200 18158
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 4080 15314 4108 17274
rect 4158 16688 4214 16697
rect 4158 16623 4160 16632
rect 4212 16623 4214 16632
rect 4160 16594 4212 16600
rect 4264 15586 4292 18702
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 4356 16522 4384 18090
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4448 17134 4476 18022
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4448 16574 4476 17070
rect 4540 16726 4568 18566
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4632 17270 4660 18022
rect 4816 17746 4844 18158
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4724 16590 4752 16934
rect 4712 16584 4764 16590
rect 4448 16546 4660 16574
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4632 16114 4660 16546
rect 4712 16526 4764 16532
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 3988 15286 4108 15314
rect 4172 15558 4292 15586
rect 3988 14550 4016 15286
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14074 4016 14350
rect 4080 14278 4108 15098
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4080 14006 4108 14214
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4080 12753 4108 13738
rect 4066 12744 4122 12753
rect 3976 12708 4028 12714
rect 4066 12679 4122 12688
rect 3976 12650 4028 12656
rect 3988 10810 4016 12650
rect 4172 12442 4200 15558
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14482 4292 14758
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 13274 4292 14418
rect 4356 14006 4384 15846
rect 4448 15706 4476 16050
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14074 4476 14758
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4448 13297 4476 13330
rect 4434 13288 4490 13297
rect 4264 13246 4384 13274
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12986 4292 13126
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4356 12918 4384 13246
rect 4434 13223 4490 13232
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4356 12714 4384 12854
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4066 12336 4122 12345
rect 4066 12271 4068 12280
rect 4120 12271 4122 12280
rect 4068 12242 4120 12248
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3882 10160 3938 10169
rect 3882 10095 3938 10104
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3330 9208 3386 9217
rect 3240 9172 3292 9178
rect 3330 9143 3386 9152
rect 3240 9114 3292 9120
rect 3252 8838 3280 9114
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3160 8622 3280 8650
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3160 6798 3188 7958
rect 3252 7886 3280 8622
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7478 3280 7686
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3056 6656 3108 6662
rect 3240 6656 3292 6662
rect 3056 6598 3108 6604
rect 3146 6624 3202 6633
rect 3240 6598 3292 6604
rect 3146 6559 3202 6568
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2976 5250 3004 6054
rect 3160 5778 3188 6559
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5409 3096 5510
rect 3054 5400 3110 5409
rect 3160 5370 3188 5714
rect 3054 5335 3110 5344
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2976 5222 3096 5250
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4282 3004 4966
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2870 4176 2926 4185
rect 2870 4111 2926 4120
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3534 2912 3878
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3068 3466 3096 5222
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3160 4622 3188 5034
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 2854 3004 3334
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2976 800 3004 2790
rect 3252 2553 3280 6598
rect 3344 2961 3372 8978
rect 3436 7970 3464 9998
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3620 9450 3648 9551
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3896 9042 3924 9386
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3988 8090 4016 10746
rect 4080 10577 4108 12242
rect 4264 11898 4292 12582
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11898 4384 12038
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4342 11112 4398 11121
rect 4342 11047 4344 11056
rect 4396 11047 4398 11056
rect 4344 11018 4396 11024
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4448 10146 4476 13126
rect 4080 10118 4476 10146
rect 4080 9897 4108 10118
rect 4160 9920 4212 9926
rect 4066 9888 4122 9897
rect 4160 9862 4212 9868
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4066 9823 4122 9832
rect 4172 9722 4200 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4172 9489 4200 9658
rect 4158 9480 4214 9489
rect 4158 9415 4214 9424
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 8673 4108 9114
rect 4448 8974 4476 9862
rect 4540 9450 4568 15982
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 12782 4660 15438
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4066 8664 4122 8673
rect 4540 8634 4568 8774
rect 4066 8599 4122 8608
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4264 8401 4292 8434
rect 4250 8392 4306 8401
rect 4250 8327 4306 8336
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4068 8016 4120 8022
rect 3436 7942 3924 7970
rect 4068 7958 4120 7964
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3436 7410 3464 7754
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3528 7290 3556 7822
rect 3436 7262 3556 7290
rect 3436 6934 3464 7262
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3330 2952 3386 2961
rect 3330 2887 3386 2896
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3238 2544 3294 2553
rect 3238 2479 3294 2488
rect 3344 800 3372 2790
rect 3436 2310 3464 6734
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6225 3832 6598
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3896 3482 3924 7942
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3988 7585 4016 7890
rect 3974 7576 4030 7585
rect 4080 7546 4108 7958
rect 3974 7511 4030 7520
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3988 6361 4016 7278
rect 4080 6934 4108 7278
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4526 6896 4582 6905
rect 4526 6831 4582 6840
rect 4540 6662 4568 6831
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3976 6248 4028 6254
rect 3974 6216 3976 6225
rect 4028 6216 4030 6225
rect 3974 6151 4030 6160
rect 4080 5914 4108 6423
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3988 5030 4016 5714
rect 4172 5370 4200 6598
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4486 4016 4966
rect 4066 4720 4122 4729
rect 4066 4655 4068 4664
rect 4120 4655 4122 4664
rect 4068 4626 4120 4632
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 3738 4016 4422
rect 4264 4298 4292 6258
rect 4540 6118 4568 6598
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4632 5914 4660 11494
rect 4724 10062 4752 14826
rect 4816 12918 4844 17546
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4908 16046 4936 16390
rect 5000 16250 5028 17478
rect 5092 16538 5120 18770
rect 5184 17882 5212 19314
rect 5736 18714 5764 22200
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 19854 7880 20334
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 7116 19417 7144 19654
rect 7944 19514 7972 19654
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7102 19408 7158 19417
rect 7102 19343 7158 19352
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6564 18834 6592 19110
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 5736 18686 5856 18714
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5538 18320 5594 18329
rect 5538 18255 5594 18264
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5184 17338 5212 17478
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5356 17128 5408 17134
rect 5354 17096 5356 17105
rect 5408 17096 5410 17105
rect 5552 17082 5580 18255
rect 5736 18057 5764 18566
rect 5828 18154 5856 18686
rect 6564 18630 6592 18770
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 5920 18222 5948 18566
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5722 18048 5778 18057
rect 5722 17983 5778 17992
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5552 17054 5672 17082
rect 5354 17031 5410 17040
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5092 16510 5212 16538
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 5092 15570 5120 16390
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5000 14618 5028 14962
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5092 14482 5120 15506
rect 5184 14793 5212 16510
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5276 14958 5304 15982
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5184 14346 5212 14554
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5276 14074 5304 14894
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5092 13734 5120 13806
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 10554 4844 12718
rect 5000 12434 5028 12786
rect 4908 12406 5028 12434
rect 4908 12102 4936 12406
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 10713 4936 12038
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4894 10704 4950 10713
rect 4894 10639 4950 10648
rect 4816 10526 4936 10554
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4816 9926 4844 10406
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4724 8498 4752 9415
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4436 4616 4488 4622
rect 4434 4584 4436 4593
rect 4488 4584 4490 4593
rect 4434 4519 4490 4528
rect 4172 4270 4292 4298
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3896 3454 4108 3482
rect 3896 3126 3924 3454
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3988 3194 4016 3334
rect 4080 3194 4108 3454
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 1737 3464 2246
rect 3422 1728 3478 1737
rect 3422 1663 3478 1672
rect 3896 1442 3924 3062
rect 4172 2774 4200 4270
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4264 3194 4292 4150
rect 4540 4060 4568 5782
rect 4632 5302 4660 5850
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 4690 4660 5102
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4758 4752 4966
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4632 4214 4660 4626
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4540 4032 4660 4060
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3602 4384 3878
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 3712 1414 3924 1442
rect 4080 2746 4200 2774
rect 3712 800 3740 1414
rect 4080 800 4108 2746
rect 4632 1442 4660 4032
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 2378 4752 3470
rect 4816 3466 4844 9862
rect 4908 8634 4936 10526
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4896 7880 4948 7886
rect 4894 7848 4896 7857
rect 4948 7848 4950 7857
rect 4894 7783 4950 7792
rect 4908 7546 4936 7783
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6458 4936 6734
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4622 4936 4966
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4816 3194 4844 3402
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5000 3126 5028 11698
rect 5092 10606 5120 13670
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 12434 5304 12582
rect 5184 12406 5304 12434
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 8430 5120 10066
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5092 6866 5120 8026
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 6118 5120 6802
rect 5184 6746 5212 12406
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5276 11694 5304 12038
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5276 9518 5304 11154
rect 5368 10742 5396 16458
rect 5460 16114 5488 16662
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 13258 5488 15098
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5552 11098 5580 14894
rect 5644 14521 5672 17054
rect 5736 16454 5764 17546
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5828 16998 5856 17274
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16794 5856 16934
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5828 16250 5856 16458
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5630 14512 5686 14521
rect 5630 14447 5686 14456
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5644 12866 5672 14282
rect 5736 14278 5764 14418
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5828 14006 5856 15914
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 12986 5764 13670
rect 5828 13326 5856 13806
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5644 12838 5764 12866
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5644 12617 5672 12650
rect 5630 12608 5686 12617
rect 5630 12543 5686 12552
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5644 11626 5672 12378
rect 5736 11830 5764 12838
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 11354 5672 11562
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5448 11076 5500 11082
rect 5552 11070 5764 11098
rect 5448 11018 5500 11024
rect 5460 10962 5488 11018
rect 5632 11008 5684 11014
rect 5460 10934 5580 10962
rect 5632 10950 5684 10956
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10130 5488 10610
rect 5552 10470 5580 10934
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7750 5304 8366
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5460 7528 5488 10066
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 8634 5580 9522
rect 5644 9042 5672 10950
rect 5736 9586 5764 11070
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5724 8968 5776 8974
rect 5644 8916 5724 8922
rect 5644 8910 5776 8916
rect 5644 8894 5764 8910
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5368 7500 5488 7528
rect 5368 6798 5396 7500
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5356 6792 5408 6798
rect 5184 6718 5304 6746
rect 5356 6734 5408 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4448 1414 4660 1442
rect 4448 800 4476 1414
rect 4816 870 4936 898
rect 4816 800 4844 870
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 4908 762 4936 870
rect 5092 762 5120 6054
rect 5184 4690 5212 6598
rect 5276 6458 5304 6718
rect 5264 6452 5316 6458
rect 5316 6412 5396 6440
rect 5264 6394 5316 6400
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5370 5304 6054
rect 5368 5914 5396 6412
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4185 5212 4422
rect 5170 4176 5226 4185
rect 5170 4111 5226 4120
rect 5184 2990 5212 4111
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5184 2650 5212 2926
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 2514 5304 3674
rect 5368 2854 5396 5850
rect 5460 5710 5488 7375
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 5914 5580 7278
rect 5644 7274 5672 8894
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 7954 5764 8774
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5644 4128 5672 6054
rect 5736 5681 5764 7686
rect 5828 6730 5856 13126
rect 5920 12442 5948 18158
rect 6012 17882 6040 18226
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6564 17678 6592 18566
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6656 17542 6684 18022
rect 6840 17626 6868 18770
rect 7300 18698 7328 19246
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7196 18624 7248 18630
rect 7116 18584 7196 18612
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6932 17746 6960 18294
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6748 17598 6868 17626
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6012 16697 6040 17478
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 5998 16688 6054 16697
rect 5998 16623 6054 16632
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6564 16250 6592 17478
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6550 15872 6606 15881
rect 6550 15807 6606 15816
rect 6564 15502 6592 15807
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6012 13530 6040 14962
rect 6564 14958 6592 15438
rect 6656 15434 6684 16458
rect 6644 15428 6696 15434
rect 6644 15370 6696 15376
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6656 14822 6684 15370
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6000 12776 6052 12782
rect 5998 12744 6000 12753
rect 6052 12744 6054 12753
rect 5998 12679 6054 12688
rect 6104 12594 6132 12786
rect 6012 12566 6132 12594
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5920 9466 5948 12174
rect 6012 10810 6040 12566
rect 6196 12238 6224 12922
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6564 11830 6592 13398
rect 6656 11898 6684 14758
rect 6748 12986 6776 17598
rect 6932 16794 6960 17682
rect 7116 17542 7144 18584
rect 7196 18566 7248 18572
rect 7300 18426 7328 18634
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7392 17610 7420 18022
rect 7470 17640 7526 17649
rect 7380 17604 7432 17610
rect 7470 17575 7526 17584
rect 7380 17546 7432 17552
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7024 16658 7052 17478
rect 7116 16726 7144 17478
rect 7392 17354 7420 17546
rect 7484 17542 7512 17575
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7392 17326 7512 17354
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16250 6868 16390
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6932 16114 6960 16526
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16182 7052 16390
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 16017 6960 16050
rect 7116 16046 7144 16458
rect 7104 16040 7156 16046
rect 6918 16008 6974 16017
rect 7104 15982 7156 15988
rect 6918 15943 6974 15952
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 13410 6868 14214
rect 6840 13382 6960 13410
rect 6932 13376 6960 13382
rect 7012 13388 7064 13394
rect 6932 13348 7012 13376
rect 7012 13330 7064 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6104 11558 6132 11630
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 9654 6040 10746
rect 6564 10538 6592 11494
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 10033 6132 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6090 10024 6146 10033
rect 6090 9959 6146 9968
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9674 6592 10202
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6472 9646 6592 9674
rect 6092 9580 6144 9586
rect 6276 9580 6328 9586
rect 6144 9540 6276 9568
rect 6092 9522 6144 9528
rect 6276 9522 6328 9528
rect 5920 9438 6040 9466
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8974 5948 9318
rect 6012 9178 6040 9438
rect 6380 9382 6408 9590
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6104 9058 6132 9318
rect 6012 9030 6132 9058
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5722 5672 5778 5681
rect 5722 5607 5778 5616
rect 5920 4146 5948 8774
rect 6012 8090 6040 9030
rect 6472 8838 6500 9646
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8362 6592 9522
rect 6656 9382 6684 10542
rect 6748 9518 6776 12650
rect 6840 12442 6868 13262
rect 7024 12850 7052 13330
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6828 12436 6880 12442
rect 7116 12434 7144 15982
rect 7208 15570 7236 16730
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14482 7236 14758
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7300 14414 7328 16934
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 16114 7420 16594
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7392 14226 7420 16050
rect 6828 12378 6880 12384
rect 7024 12406 7144 12434
rect 7208 14198 7420 14226
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 11762 6868 12242
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6932 11218 6960 12038
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6840 9042 6868 11154
rect 6932 11121 6960 11154
rect 6918 11112 6974 11121
rect 6918 11047 6974 11056
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6564 8022 6592 8298
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6012 7546 6040 7686
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6012 6254 6040 6802
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6012 5846 6040 6190
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6012 5166 6040 5782
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6472 5681 6500 5714
rect 6458 5672 6514 5681
rect 6458 5607 6514 5616
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6564 4622 6592 7686
rect 6656 5409 6684 8774
rect 6840 7313 6868 8978
rect 6932 8906 6960 9318
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 7024 8514 7052 12406
rect 7104 12096 7156 12102
rect 7102 12064 7104 12073
rect 7156 12064 7158 12073
rect 7102 11999 7158 12008
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7116 10266 7144 11834
rect 7208 10690 7236 14198
rect 7484 13802 7512 17326
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7576 13433 7604 19110
rect 8036 18426 8064 19246
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8312 18426 8340 18702
rect 8496 18426 8524 19858
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8496 18222 8524 18362
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17218 8340 18090
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17338 8432 17478
rect 8496 17338 8524 18022
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8312 17190 8524 17218
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 7746 16552 7802 16561
rect 7746 16487 7802 16496
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7668 15910 7696 16186
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7562 13424 7618 13433
rect 7562 13359 7618 13368
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11082 7328 12582
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7392 10826 7420 12922
rect 7484 11898 7512 13126
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7576 12102 7604 12242
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7392 10798 7512 10826
rect 7208 10662 7420 10690
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6932 8498 7052 8514
rect 6920 8492 7052 8498
rect 6972 8486 7052 8492
rect 6920 8434 6972 8440
rect 7024 8022 7052 8486
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7116 7954 7144 8774
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6826 7304 6882 7313
rect 6826 7239 6882 7248
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 6882 6960 7142
rect 7024 7002 7052 7686
rect 7208 7410 7236 10406
rect 7300 10266 7328 10542
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7300 8430 7328 9114
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7478 7328 7890
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7392 7188 7420 10662
rect 7300 7160 7420 7188
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6828 6860 6880 6866
rect 6932 6854 7052 6882
rect 6828 6802 6880 6808
rect 6840 6118 6868 6802
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6322 6960 6734
rect 7024 6662 7052 6854
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6390 7052 6598
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7116 6254 7144 6734
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6642 5400 6698 5409
rect 6642 5335 6698 5344
rect 6748 5284 6776 5510
rect 6840 5370 6868 6054
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6656 5256 6776 5284
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 5460 4100 5672 4128
rect 5908 4140 5960 4146
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 4908 734 5120 762
rect 5170 0 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 4100
rect 5908 4082 5960 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5724 3664 5776 3670
rect 5538 3632 5594 3641
rect 5724 3606 5776 3612
rect 5538 3567 5540 3576
rect 5592 3567 5594 3576
rect 5540 3538 5592 3544
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5552 2446 5580 3402
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5552 800 5580 2382
rect 5644 2378 5672 2858
rect 5736 2854 5764 3606
rect 5828 3097 5856 4014
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3466 5948 3878
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3194 5948 3402
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5814 3088 5870 3097
rect 5814 3023 5870 3032
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 6012 2774 6040 3946
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 5920 2746 6040 2774
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5920 800 5948 2746
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6288 870 6408 898
rect 6288 800 6316 870
rect 5276 734 5488 762
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6380 762 6408 870
rect 6564 762 6592 4082
rect 6656 800 6684 5256
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7116 4826 7144 5170
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6748 3233 6776 3606
rect 7024 3534 7052 4014
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7010 3360 7066 3369
rect 6734 3224 6790 3233
rect 6734 3159 6790 3168
rect 6932 3126 6960 3334
rect 7010 3295 7066 3304
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6918 2544 6974 2553
rect 6918 2479 6974 2488
rect 6932 2446 6960 2479
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7024 800 7052 3295
rect 7208 2446 7236 4490
rect 7300 4078 7328 7160
rect 7484 6798 7512 10798
rect 7576 7206 7604 12038
rect 7668 11898 7696 15506
rect 7760 15366 7788 16487
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 14770 7788 15302
rect 7852 14958 7880 17002
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8036 16697 8064 16934
rect 8404 16794 8432 17002
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8300 16720 8352 16726
rect 8022 16688 8078 16697
rect 7932 16652 7984 16658
rect 8300 16662 8352 16668
rect 8022 16623 8078 16632
rect 7932 16594 7984 16600
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7760 14742 7880 14770
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12782 7788 13126
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7852 12628 7880 14742
rect 7760 12600 7880 12628
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 10849 7788 12600
rect 7944 11830 7972 16594
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8036 15706 8064 15982
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8128 15586 8156 16118
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8036 15558 8156 15586
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7944 11150 7972 11630
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7746 10840 7802 10849
rect 7746 10775 7802 10784
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7668 8838 7696 10066
rect 7760 10062 7788 10542
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7654 8120 7710 8129
rect 7654 8055 7656 8064
rect 7708 8055 7710 8064
rect 7656 8026 7708 8032
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6934 7604 7142
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7760 6390 7788 9998
rect 7852 8634 7880 10950
rect 7930 10840 7986 10849
rect 7930 10775 7986 10784
rect 7944 10033 7972 10775
rect 7930 10024 7986 10033
rect 8036 9994 8064 15558
rect 8220 15366 8248 15846
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8206 14784 8262 14793
rect 8206 14719 8262 14728
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8128 13190 8156 13466
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12918 8156 13126
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 8128 12238 8156 12854
rect 8220 12646 8248 14719
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8208 12096 8260 12102
rect 8206 12064 8208 12073
rect 8260 12064 8262 12073
rect 8206 11999 8262 12008
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7930 9959 7986 9968
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 6662 7880 7142
rect 8036 6866 8064 8978
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7392 5914 7420 6190
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5778 7512 6190
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3602 7328 3878
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7300 1834 7328 3538
rect 7484 2774 7512 5714
rect 7576 5642 7604 6258
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7760 5574 7788 6326
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7392 2746 7512 2774
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 7392 800 7420 2746
rect 7576 2514 7604 3470
rect 7668 3058 7696 5102
rect 7852 4486 7880 6598
rect 8128 5710 8156 11494
rect 8220 9654 8248 11766
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8206 8936 8262 8945
rect 8206 8871 8262 8880
rect 8220 8634 8248 8871
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8220 7546 8248 7890
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8022 5536 8078 5545
rect 8022 5471 8078 5480
rect 8036 4622 8064 5471
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7760 2961 7788 3334
rect 7746 2952 7802 2961
rect 7746 2887 7802 2896
rect 7852 2774 7880 4422
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7944 4049 7972 4218
rect 7930 4040 7986 4049
rect 7930 3975 7986 3984
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8128 3534 8156 3674
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7760 2746 7880 2774
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7760 800 7788 2746
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 7852 1970 7880 2246
rect 8036 2106 8064 2246
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 8128 800 8156 3062
rect 8220 3058 8248 7278
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8312 2774 8340 16662
rect 8404 14414 8432 16730
rect 8496 15570 8524 17190
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 5234 8432 14214
rect 8496 12434 8524 15030
rect 8588 12986 8616 19314
rect 9876 19310 9904 19790
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 9968 19417 9996 19654
rect 10428 19514 10456 19654
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9954 19408 10010 19417
rect 9954 19343 10010 19352
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8956 18290 8984 18770
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8680 17338 8708 18226
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8772 17542 8800 17818
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8680 16182 8708 17070
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8772 15994 8800 16662
rect 8680 15966 8800 15994
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8680 12434 8708 15966
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8772 15162 8800 15506
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 9232 15026 9260 15438
rect 9324 15434 9352 19246
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9416 17882 9444 18158
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9508 17746 9536 18158
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 17202 9444 17546
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9416 16726 9444 17138
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 14006 8800 14214
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8956 13938 8984 14350
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8496 12406 8616 12434
rect 8680 12406 8984 12434
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11082 8524 11494
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8588 10826 8616 12406
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8680 11830 8708 12310
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8680 11150 8708 11766
rect 8956 11540 8984 12406
rect 9140 12374 9168 14486
rect 9232 14482 9260 14962
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9232 13938 9260 14418
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9232 13394 9260 13874
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 8956 11512 9168 11540
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8588 10798 8708 10826
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 9926 8616 10610
rect 8680 10538 8708 10798
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8496 8906 8524 9386
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 8294 8524 8434
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 6730 8524 7686
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8588 6322 8616 9862
rect 8680 8974 8708 10474
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9140 9738 9168 11512
rect 9048 9710 9168 9738
rect 9048 9489 9076 9710
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9034 9480 9090 9489
rect 9034 9415 9090 9424
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8668 8968 8720 8974
rect 8720 8916 8800 8922
rect 8668 8910 8800 8916
rect 8680 8894 8800 8910
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 7818 8708 8502
rect 8772 8294 8800 8894
rect 9048 8362 9076 8978
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8680 6202 8708 7754
rect 9140 7206 9168 9590
rect 9232 9330 9260 13194
rect 9324 12986 9352 14282
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 10810 9352 12582
rect 9416 11286 9444 15846
rect 9508 14346 9536 17682
rect 9692 17542 9720 18566
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17610 9812 17818
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9600 17270 9628 17478
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9496 13932 9548 13938
rect 9600 13920 9628 17070
rect 9548 13892 9628 13920
rect 9496 13874 9548 13880
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9324 9994 9352 10746
rect 9416 10266 9444 11222
rect 9508 11150 9536 11834
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9416 9654 9444 10202
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9232 9302 9444 9330
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 8294 9260 8366
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9324 7886 9352 9046
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9232 7410 9260 7822
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9232 7002 9260 7346
rect 9310 7304 9366 7313
rect 9310 7239 9366 7248
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 8852 6384 8904 6390
rect 8850 6352 8852 6361
rect 8904 6352 8906 6361
rect 8850 6287 8906 6296
rect 8852 6248 8904 6254
rect 8588 6174 8708 6202
rect 8758 6216 8814 6225
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8588 4146 8616 6174
rect 8814 6196 8852 6202
rect 8814 6190 8904 6196
rect 8942 6216 8998 6225
rect 8814 6174 8892 6190
rect 8758 6151 8814 6160
rect 8942 6151 8944 6160
rect 8996 6151 8998 6160
rect 8944 6122 8996 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8496 3942 8524 4082
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8588 3398 8616 4082
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8312 2746 8524 2774
rect 8496 800 8524 2746
rect 8588 2514 8616 3334
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8680 2446 8708 5578
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9140 4282 9168 6598
rect 9324 5846 9352 7239
rect 9416 6662 9444 9302
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9508 7970 9536 8502
rect 9600 8090 9628 13892
rect 9692 12889 9720 17478
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9784 15026 9812 16186
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9678 12880 9734 12889
rect 9678 12815 9734 12824
rect 9784 12730 9812 14554
rect 9876 13258 9904 19246
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18290 9996 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9968 17338 9996 18226
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 14278 10088 18362
rect 10152 18057 10180 19246
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18086 10364 18634
rect 10324 18080 10376 18086
rect 10138 18048 10194 18057
rect 10324 18022 10376 18028
rect 10138 17983 10194 17992
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16250 10180 16390
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10152 14414 10180 16186
rect 10244 15706 10272 17682
rect 10336 17610 10364 18022
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10428 17338 10456 17478
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9968 13138 9996 14214
rect 10060 13938 10088 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9692 12702 9812 12730
rect 9876 13110 9996 13138
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9692 12345 9720 12702
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10470 9720 11018
rect 9680 10464 9732 10470
rect 9732 10412 9812 10418
rect 9680 10406 9812 10412
rect 9692 10390 9812 10406
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9518 9720 9998
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9784 9330 9812 10390
rect 9692 9302 9812 9330
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9508 7942 9628 7970
rect 9600 6905 9628 7942
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9600 6361 9628 6394
rect 9586 6352 9642 6361
rect 9404 6316 9456 6322
rect 9586 6287 9642 6296
rect 9404 6258 9456 6264
rect 9416 6118 9444 6258
rect 9692 6186 9720 9302
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9784 8906 9812 9114
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9876 7993 9904 13110
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9968 11354 9996 12922
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9968 10266 9996 10678
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10060 9654 10088 13126
rect 10152 12628 10180 13670
rect 10244 12918 10272 15642
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10232 12640 10284 12646
rect 10152 12600 10232 12628
rect 10232 12582 10284 12588
rect 10138 11792 10194 11801
rect 10138 11727 10140 11736
rect 10192 11727 10194 11736
rect 10140 11698 10192 11704
rect 10244 10554 10272 12582
rect 10336 12170 10364 14758
rect 10428 12986 10456 14962
rect 10520 14414 10548 19858
rect 12360 19854 12388 20198
rect 13740 20058 13768 20470
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14384 20058 14412 20402
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 11072 19718 11100 19790
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11060 19712 11112 19718
rect 11058 19680 11060 19689
rect 11704 19712 11756 19718
rect 11112 19680 11114 19689
rect 11704 19654 11756 19660
rect 11058 19615 11114 19624
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11610 18864 11666 18873
rect 10968 18828 11020 18834
rect 11610 18799 11666 18808
rect 10968 18770 11020 18776
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 17338 10640 17546
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10612 16114 10640 17274
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15570 10640 16050
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 13530 10548 14350
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10506 13288 10562 13297
rect 10506 13223 10562 13232
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10414 12744 10470 12753
rect 10414 12679 10470 12688
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10152 10526 10272 10554
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 8974 9996 9318
rect 10060 9178 10088 9590
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9784 6798 9812 7210
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 9324 5574 9352 5607
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4690 9260 5306
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9416 4570 9444 6054
rect 9692 5681 9720 6122
rect 9678 5672 9734 5681
rect 10060 5642 10088 7142
rect 9678 5607 9734 5616
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9232 4542 9444 4570
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8942 4176 8998 4185
rect 8942 4111 8944 4120
rect 8996 4111 8998 4120
rect 8944 4082 8996 4088
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8864 3466 8892 3674
rect 9232 3516 9260 4542
rect 9402 4176 9458 4185
rect 9402 4111 9458 4120
rect 9310 4040 9366 4049
rect 9310 3975 9312 3984
rect 9364 3975 9366 3984
rect 9312 3946 9364 3952
rect 9416 3942 9444 4111
rect 9588 4072 9640 4078
rect 9586 4040 9588 4049
rect 9640 4040 9642 4049
rect 9784 4010 9812 4694
rect 9586 3975 9642 3984
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9404 3936 9456 3942
rect 9456 3884 9536 3890
rect 9404 3878 9536 3884
rect 9416 3862 9536 3878
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 8942 3496 8998 3505
rect 8852 3460 8904 3466
rect 8942 3431 8998 3440
rect 9140 3488 9260 3516
rect 8852 3402 8904 3408
rect 8956 3398 8984 3431
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9048 2836 9076 3334
rect 9140 2938 9168 3488
rect 9218 3360 9274 3369
rect 9218 3295 9274 3304
rect 9232 3058 9260 3295
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9140 2910 9260 2938
rect 9048 2808 9168 2836
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9140 2446 9168 2808
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 800 8892 2246
rect 9232 800 9260 2910
rect 9324 1426 9352 3606
rect 9508 3398 9536 3862
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9508 2378 9536 3062
rect 9784 3058 9812 3946
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9876 2938 9904 3878
rect 9692 2910 9904 2938
rect 9692 2854 9720 2910
rect 9680 2848 9732 2854
rect 9772 2848 9824 2854
rect 9680 2790 9732 2796
rect 9770 2816 9772 2825
rect 9824 2816 9826 2825
rect 9770 2751 9826 2760
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9588 1692 9640 1698
rect 9588 1634 9640 1640
rect 9312 1420 9364 1426
rect 9312 1362 9364 1368
rect 9600 800 9628 1634
rect 9968 800 9996 5578
rect 10152 5234 10180 10526
rect 10336 10266 10364 12106
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10428 9654 10456 12679
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10520 9382 10548 13223
rect 10704 11082 10732 17682
rect 10796 16153 10824 18022
rect 10980 16697 11008 18770
rect 11624 18766 11652 18799
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11072 18329 11100 18566
rect 11058 18320 11114 18329
rect 11058 18255 11114 18264
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10966 16688 11022 16697
rect 10966 16623 10968 16632
rect 11020 16623 11022 16632
rect 10968 16594 11020 16600
rect 10782 16144 10838 16153
rect 10782 16079 10838 16088
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15502 10824 15846
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10888 14618 10916 14826
rect 10980 14618 11008 15370
rect 11072 14822 11100 17750
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16726 11192 16934
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11256 16590 11284 18566
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11716 15638 11744 18634
rect 11900 18222 11928 19722
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12084 18630 12112 18838
rect 12360 18766 12388 19246
rect 12452 18902 12480 19858
rect 12636 19514 12664 19926
rect 13740 19922 13768 19994
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12348 18760 12400 18766
rect 12636 18737 12664 18770
rect 12348 18702 12400 18708
rect 12622 18728 12678 18737
rect 12622 18663 12678 18672
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18426 12848 18566
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 13556 18290 13584 18906
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11900 17134 11928 18158
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11256 14550 11284 14758
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11716 13870 11744 14758
rect 11808 14278 11836 17070
rect 11900 16658 11928 17070
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13938 11836 14214
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11704 13864 11756 13870
rect 11900 13818 11928 16594
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11704 13806 11756 13812
rect 11716 13190 11744 13806
rect 11808 13790 11928 13818
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12986 11744 13126
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 10888 12850 10916 12922
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10888 12306 10916 12786
rect 11808 12442 11836 13790
rect 11992 13682 12020 14486
rect 11900 13654 12020 13682
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10888 11762 10916 12242
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11716 11778 11744 11834
rect 11900 11830 11928 13654
rect 11888 11824 11940 11830
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10888 11354 10916 11698
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10704 10577 10732 10610
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8294 10272 8910
rect 10428 8906 10456 8978
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10322 8256 10378 8265
rect 10244 7886 10272 8230
rect 10322 8191 10378 8200
rect 10232 7880 10284 7886
rect 10336 7857 10364 8191
rect 10232 7822 10284 7828
rect 10322 7848 10378 7857
rect 10322 7783 10378 7792
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 2446 10088 4422
rect 10152 3602 10180 5170
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10152 2446 10180 2926
rect 10244 2825 10272 5510
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 1902 10180 2246
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10336 800 10364 7783
rect 10428 4758 10456 8842
rect 10612 8294 10640 9959
rect 10796 9926 10824 11222
rect 10888 10606 10916 11290
rect 10876 10600 10928 10606
rect 10928 10560 11008 10588
rect 10876 10542 10928 10548
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10796 7546 10824 9862
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10692 7472 10744 7478
rect 10888 7426 10916 9590
rect 10980 8974 11008 10560
rect 11164 9994 11192 11766
rect 11624 11626 11652 11766
rect 11716 11750 11836 11778
rect 11888 11766 11940 11772
rect 11808 11642 11836 11750
rect 11612 11620 11664 11626
rect 11808 11614 11928 11642
rect 11612 11562 11664 11568
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11164 9722 11192 9930
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11624 8974 11652 9386
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11808 8838 11836 8978
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11152 7880 11204 7886
rect 10692 7414 10744 7420
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10520 1698 10548 6666
rect 10612 4282 10640 7414
rect 10704 4690 10732 7414
rect 10796 7398 10916 7426
rect 10980 7840 11152 7868
rect 10796 5030 10824 7398
rect 10980 7313 11008 7840
rect 11152 7822 11204 7828
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 10966 7304 11022 7313
rect 10966 7239 11022 7248
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11072 6798 11100 7142
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6662 11100 6734
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11058 5400 11114 5409
rect 11058 5335 11114 5344
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4729 10824 4966
rect 10782 4720 10838 4729
rect 10692 4684 10744 4690
rect 10782 4655 10838 4664
rect 10692 4626 10744 4632
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10612 3738 10640 4218
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10690 3904 10746 3913
rect 10690 3839 10746 3848
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10508 1692 10560 1698
rect 10508 1634 10560 1640
rect 10704 800 10732 3839
rect 10888 3738 10916 4150
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 2038 10916 2246
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 11072 800 11100 5335
rect 11164 4554 11192 7142
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 5574 11284 6666
rect 11716 6662 11744 7686
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11716 6254 11744 6598
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11716 5574 11744 6190
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11716 5302 11744 5510
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4010 11192 4490
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11150 3904 11206 3913
rect 11150 3839 11206 3848
rect 11164 3058 11192 3839
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2650 11192 2994
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2446 11284 5034
rect 11716 5030 11744 5238
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4622 11744 4966
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11716 4146 11744 4558
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11348 3942 11376 4082
rect 11336 3936 11388 3942
rect 11334 3904 11336 3913
rect 11388 3904 11390 3913
rect 11334 3839 11390 3848
rect 11348 3813 11376 3839
rect 11808 3466 11836 8298
rect 11612 3460 11664 3466
rect 11796 3460 11848 3466
rect 11664 3420 11744 3448
rect 11612 3402 11664 3408
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11716 3058 11744 3420
rect 11796 3402 11848 3408
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 6380 734 6592 762
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 2994
rect 11900 2774 11928 11614
rect 12084 11218 12112 16186
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12442 12296 13194
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10169 12204 10678
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12360 9674 12388 17750
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12820 14074 12848 16594
rect 13004 16590 13032 16934
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12912 13870 12940 14214
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 10674 12480 12582
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12268 9646 12388 9674
rect 12268 8945 12296 9646
rect 12452 9586 12480 9862
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 12164 8288 12216 8294
rect 13096 8265 13124 15846
rect 13280 15502 13308 16934
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13280 14822 13308 15098
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 13188 12374 13216 12679
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11898 13216 12310
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13280 9178 13308 12106
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 8430 13308 8842
rect 13372 8430 13400 16390
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13464 15706 13492 16186
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13556 15473 13584 17478
rect 13542 15464 13598 15473
rect 13542 15399 13598 15408
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13464 14550 13492 14826
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13556 14414 13584 14962
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 14278 13584 14350
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13648 12434 13676 19790
rect 14568 19718 14596 19994
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 16250 13768 18226
rect 13832 17270 13860 18362
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 14292 17338 14320 17546
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 14292 16998 14320 17274
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13740 14618 13768 16050
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13556 12406 13676 12434
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11218 13492 11698
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12164 8230 12216 8236
rect 13082 8256 13138 8265
rect 12176 8090 12204 8230
rect 13082 8191 13138 8200
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 5914 12020 6734
rect 13464 6458 13492 7346
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12176 4826 12204 6258
rect 13464 6118 13492 6394
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5098 12480 5578
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12176 4214 12204 4490
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3670 12112 3878
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12452 3466 12480 5034
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12440 2984 12492 2990
rect 12544 2972 12572 3674
rect 12636 3534 12664 4694
rect 13082 4176 13138 4185
rect 13464 4146 13492 5714
rect 13082 4111 13084 4120
rect 13136 4111 13138 4120
rect 13452 4140 13504 4146
rect 13084 4082 13136 4088
rect 13452 4082 13504 4088
rect 13266 3632 13322 3641
rect 13266 3567 13322 3576
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 13280 3194 13308 3567
rect 13556 3194 13584 12406
rect 13832 12238 13860 12718
rect 13924 12646 13952 12922
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11830 13860 12174
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 14278 11656 14334 11665
rect 14278 11591 14334 11600
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13832 10606 13860 11086
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13832 10062 13860 10542
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14292 9178 14320 11591
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 13740 8974 13768 9114
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7206 13676 8230
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 6798 13676 7142
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6118 13676 6734
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5250 13676 6054
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5386 13860 5510
rect 13740 5370 13860 5386
rect 13728 5364 13860 5370
rect 13780 5358 13860 5364
rect 13728 5306 13780 5312
rect 13648 5234 13768 5250
rect 13648 5228 13780 5234
rect 13648 5222 13728 5228
rect 13728 5170 13780 5176
rect 13740 4690 13768 5170
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13740 3942 13768 4626
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3652 13768 3878
rect 13832 3777 13860 5358
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13818 3768 13874 3777
rect 13945 3771 14253 3780
rect 13818 3703 13874 3712
rect 13740 3624 13860 3652
rect 13832 3534 13860 3624
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12492 2944 12572 2972
rect 12440 2926 12492 2932
rect 11808 2746 11928 2774
rect 11808 800 11836 2746
rect 12452 2650 12480 2926
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12176 800 12204 2450
rect 12532 2100 12584 2106
rect 12532 2042 12584 2048
rect 12544 800 12572 2042
rect 12912 800 12940 3062
rect 14292 3058 14320 8366
rect 14384 3738 14412 19382
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14476 18970 14504 19314
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 15502 14504 18158
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 13734 14504 14214
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13530 14504 13670
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14476 12442 14504 12786
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 10266 14504 12378
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 9722 14504 10202
rect 14568 10198 14596 13398
rect 14660 11121 14688 18906
rect 14752 18170 14780 19858
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19514 14872 19790
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15396 19378 15424 19722
rect 16040 19514 16068 19858
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18766 15240 19110
rect 15016 18760 15068 18766
rect 15200 18760 15252 18766
rect 15068 18720 15148 18748
rect 15016 18702 15068 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14752 18142 14872 18170
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14646 11112 14702 11121
rect 14646 11047 14702 11056
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14476 7818 14504 8434
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 3942 14504 5578
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14476 3097 14504 3878
rect 14462 3088 14518 3097
rect 14280 3052 14332 3058
rect 14752 3058 14780 18022
rect 14844 15162 14872 18142
rect 15028 16250 15056 18566
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14844 11830 14872 15098
rect 15120 12434 15148 18720
rect 15200 18702 15252 18708
rect 15212 17882 15240 18702
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15396 18426 15424 18566
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15304 17338 15332 18226
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15488 17218 15516 19246
rect 16040 18714 16068 19450
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16500 18970 16528 19178
rect 16960 18970 16988 19654
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16946 18864 17002 18873
rect 16120 18828 16172 18834
rect 17144 18834 17172 19450
rect 17236 19174 17264 22200
rect 19522 21312 19578 21321
rect 19522 21247 19578 21256
rect 18050 20496 18106 20505
rect 18050 20431 18106 20440
rect 18236 20460 18288 20466
rect 17408 20256 17460 20262
rect 17408 20198 17460 20204
rect 17420 19854 17448 20198
rect 18064 20058 18092 20431
rect 18236 20402 18288 20408
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 20262 18184 20334
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17960 19984 18012 19990
rect 17958 19952 17960 19961
rect 18012 19952 18014 19961
rect 17684 19916 17736 19922
rect 17958 19887 18014 19896
rect 17684 19858 17736 19864
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17512 19417 17540 19654
rect 17604 19514 17632 19654
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17498 19408 17554 19417
rect 17498 19343 17554 19352
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 16946 18799 17002 18808
rect 17132 18828 17184 18834
rect 16120 18770 16172 18776
rect 15948 18686 16068 18714
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15028 12406 15148 12434
rect 15212 17190 15516 17218
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14936 11694 14964 12174
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 10554 14964 10610
rect 15028 10554 15056 12406
rect 15212 10810 15240 17190
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15290 16688 15346 16697
rect 15290 16623 15346 16632
rect 15304 14074 15332 16623
rect 15396 15366 15424 17002
rect 15764 16794 15792 17478
rect 15856 17338 15884 17614
rect 15844 17332 15896 17338
rect 15844 17274 15896 17280
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15488 15094 15516 16594
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15476 15088 15528 15094
rect 15382 15056 15438 15065
rect 15476 15030 15528 15036
rect 15382 14991 15438 15000
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12170 15332 12582
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 14936 10526 15056 10554
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8566 14964 8774
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 15028 7206 15056 10526
rect 15396 9602 15424 14991
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14618 15516 14894
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15396 9574 15516 9602
rect 15580 9586 15608 16458
rect 15672 14618 15700 16730
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15764 14414 15792 14758
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 13870 15792 14350
rect 15856 14346 15884 15302
rect 15948 15162 15976 18686
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 16522 16068 18566
rect 16132 17066 16160 18770
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18086 16252 18702
rect 16960 18698 16988 18799
rect 17132 18770 17184 18776
rect 17236 18748 17264 19110
rect 17406 18864 17462 18873
rect 17406 18799 17462 18808
rect 17236 18720 17356 18748
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15672 12374 15700 12854
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15764 12238 15792 12786
rect 15948 12434 15976 15098
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 14074 16068 14350
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16040 13326 16068 13806
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16040 12986 16068 13262
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15856 12406 15976 12434
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10470 15792 10950
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10062 15792 10406
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 8974 15424 9454
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15120 8294 15148 8570
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7274 15332 7890
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 3602 15056 7142
rect 15488 6458 15516 9574
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15856 9058 15884 12406
rect 16132 11642 16160 15846
rect 16224 14958 16252 18022
rect 16316 15910 16344 18022
rect 16408 17814 16436 18634
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16486 18184 16542 18193
rect 16960 18154 16988 18634
rect 16486 18119 16542 18128
rect 16948 18148 17000 18154
rect 16500 17882 16528 18119
rect 16948 18090 17000 18096
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16408 16658 16436 17614
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16868 16538 16896 17274
rect 16960 17202 16988 18090
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16658 16988 16934
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16868 16510 16988 16538
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 16250 16436 16390
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16960 15706 16988 16510
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16316 11898 16344 15642
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15162 16988 15438
rect 17052 15434 17080 16594
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16408 13258 16436 14554
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16960 13410 16988 14758
rect 17052 13530 17080 15370
rect 17236 15026 17264 15642
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17236 14090 17264 14962
rect 17328 14822 17356 18720
rect 17420 18358 17448 18799
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18358 17540 18566
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17420 14618 17448 18158
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17236 14062 17356 14090
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16960 13382 17080 13410
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16132 11614 16344 11642
rect 16316 11558 16344 11614
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15764 9030 15884 9058
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15672 7886 15700 8842
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15580 6338 15608 7142
rect 15764 6662 15792 9030
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8430 15884 8910
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15856 8294 15884 8366
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7954 15884 8230
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6338 15792 6598
rect 15948 6474 15976 9454
rect 16040 8974 16068 10746
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 15488 6310 15608 6338
rect 15672 6310 15792 6338
rect 15856 6446 15976 6474
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15120 3482 15148 3538
rect 15028 3454 15148 3482
rect 14462 3023 14518 3032
rect 14740 3052 14792 3058
rect 14280 2994 14332 3000
rect 14740 2994 14792 3000
rect 13176 2984 13228 2990
rect 14188 2984 14240 2990
rect 13176 2926 13228 2932
rect 13818 2952 13874 2961
rect 13188 2650 13216 2926
rect 14240 2932 14320 2938
rect 14188 2926 14320 2932
rect 14200 2910 14320 2926
rect 13818 2887 13874 2896
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13280 2106 13308 2518
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13280 800 13308 1906
rect 13556 1834 13584 2450
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13832 1442 13860 2887
rect 14292 2854 14320 2910
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14292 2650 14320 2790
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 13636 1420 13688 1426
rect 13832 1414 14044 1442
rect 13636 1362 13688 1368
rect 13648 800 13676 1362
rect 14016 800 14044 1414
rect 14384 800 14412 2382
rect 14752 800 14780 2858
rect 15028 2378 15056 3454
rect 15212 2990 15240 4422
rect 15304 4282 15332 5306
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15488 5250 15516 6310
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 5370 15608 5646
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15396 4321 15424 5238
rect 15488 5222 15608 5250
rect 15580 5098 15608 5222
rect 15568 5092 15620 5098
rect 15568 5034 15620 5040
rect 15382 4312 15438 4321
rect 15292 4276 15344 4282
rect 15382 4247 15438 4256
rect 15292 4218 15344 4224
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15304 3942 15332 4082
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15580 3670 15608 5034
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15120 2446 15148 2926
rect 15212 2650 15240 2926
rect 15672 2922 15700 6310
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5574 15792 6190
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15764 2774 15792 3062
rect 15672 2746 15792 2774
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15672 2514 15700 2746
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 15856 2446 15884 6446
rect 15936 6384 15988 6390
rect 15934 6352 15936 6361
rect 15988 6352 15990 6361
rect 15934 6287 15990 6296
rect 16040 3126 16068 6666
rect 16132 6322 16160 7822
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16132 4826 16160 6258
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4010 16252 9318
rect 16316 7274 16344 11494
rect 16684 11150 16712 11494
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9586 16436 10066
rect 16960 9994 16988 12038
rect 17052 10266 17080 13382
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 11370 17172 13126
rect 17236 12102 17264 13874
rect 17328 13190 17356 14062
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17144 11354 17264 11370
rect 17144 11348 17276 11354
rect 17144 11342 17224 11348
rect 17224 11290 17276 11296
rect 17420 11082 17448 14554
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 17052 9654 17080 10202
rect 17144 9926 17172 10610
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17052 8838 17080 8978
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 17144 8634 17172 9862
rect 17512 9674 17540 18294
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17604 13530 17632 13874
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17604 12850 17632 13466
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17604 12442 17632 12786
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17328 9646 17540 9674
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16316 5166 16344 7210
rect 16408 7206 16436 8230
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16948 6248 17000 6254
rect 17052 6225 17080 6258
rect 16948 6190 17000 6196
rect 17038 6216 17094 6225
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16408 4010 16436 6190
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16578 5264 16634 5273
rect 16578 5199 16580 5208
rect 16632 5199 16634 5208
rect 16580 5170 16632 5176
rect 16868 4622 16896 5306
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16592 3534 16620 3674
rect 16672 3664 16724 3670
rect 16670 3632 16672 3641
rect 16724 3632 16726 3641
rect 16670 3567 16726 3576
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3194 16344 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16960 3194 16988 6190
rect 17038 6151 17094 6160
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15120 800 15148 1838
rect 11532 734 11744 762
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15212 762 15240 2246
rect 15844 2032 15896 2038
rect 15844 1974 15896 1980
rect 15396 870 15516 898
rect 15396 762 15424 870
rect 15488 800 15516 870
rect 15856 800 15884 1974
rect 16224 800 16252 2858
rect 17144 2446 17172 6598
rect 17236 5642 17264 8774
rect 17328 7970 17356 9646
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17420 8294 17448 8774
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17328 7942 17540 7970
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 6798 17356 7686
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17420 6458 17448 7822
rect 17512 7449 17540 7942
rect 17604 7546 17632 12106
rect 17696 10810 17724 19858
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 18970 17816 19246
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17774 18320 17830 18329
rect 17774 18255 17830 18264
rect 17788 17882 17816 18255
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17498 7440 17554 7449
rect 17498 7375 17554 7384
rect 17696 6633 17724 9114
rect 17788 7970 17816 15982
rect 17880 15178 17908 19110
rect 18156 18834 18184 20198
rect 18248 19922 18276 20402
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18524 19446 18552 20198
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 19514 18736 19654
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18524 18970 18552 19382
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 18064 17678 18092 18634
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18052 17264 18104 17270
rect 18050 17232 18052 17241
rect 18104 17232 18106 17241
rect 18050 17167 18106 17176
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16697 18000 17002
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 18064 16538 18092 17070
rect 17972 16522 18092 16538
rect 17960 16516 18092 16522
rect 18012 16510 18092 16516
rect 17960 16458 18012 16464
rect 17972 15858 18000 16458
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 15978 18092 16390
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 17972 15830 18092 15858
rect 17880 15150 18000 15178
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11150 17908 11630
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10674 17908 11086
rect 17972 10826 18000 15150
rect 18064 12345 18092 15830
rect 18156 13190 18184 18770
rect 18236 18760 18288 18766
rect 18234 18728 18236 18737
rect 18288 18728 18290 18737
rect 18234 18663 18290 18672
rect 18340 18290 18368 18906
rect 18524 18426 18552 18906
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18248 17746 18276 18022
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18234 16144 18290 16153
rect 18234 16079 18290 16088
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18050 12336 18106 12345
rect 18050 12271 18106 12280
rect 18156 12102 18184 13126
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18248 11914 18276 16079
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18340 14822 18368 15302
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14278 18368 14758
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 13938 18368 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18156 11886 18276 11914
rect 18050 11792 18106 11801
rect 18050 11727 18052 11736
rect 18104 11727 18106 11736
rect 18052 11698 18104 11704
rect 17972 10798 18092 10826
rect 18064 10742 18092 10798
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 10062 17908 10610
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17868 10056 17920 10062
rect 17972 10033 18000 10202
rect 17868 9998 17920 10004
rect 17958 10024 18014 10033
rect 17958 9959 18014 9968
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17868 9104 17920 9110
rect 17972 9081 18000 9522
rect 17868 9046 17920 9052
rect 17958 9072 18014 9081
rect 17880 8634 17908 9046
rect 17958 9007 18014 9016
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 8090 18000 8842
rect 18064 8106 18092 10678
rect 18156 8537 18184 11886
rect 18142 8528 18198 8537
rect 18142 8463 18198 8472
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 17960 8084 18012 8090
rect 18064 8078 18184 8106
rect 17960 8026 18012 8032
rect 17788 7942 17908 7970
rect 17774 7848 17830 7857
rect 17774 7783 17830 7792
rect 17682 6624 17738 6633
rect 17682 6559 17738 6568
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17788 6338 17816 7783
rect 17604 6310 17816 6338
rect 17500 5704 17552 5710
rect 17314 5672 17370 5681
rect 17224 5636 17276 5642
rect 17500 5646 17552 5652
rect 17314 5607 17370 5616
rect 17224 5578 17276 5584
rect 17328 5234 17356 5607
rect 17512 5370 17540 5646
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4826 17356 5170
rect 17316 4820 17368 4826
rect 17236 4780 17316 4808
rect 17236 2990 17264 4780
rect 17316 4762 17368 4768
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17328 3602 17356 4082
rect 17604 3738 17632 6310
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17696 4078 17724 5578
rect 17788 4185 17816 6122
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17880 3738 17908 7942
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18064 7449 18092 7890
rect 18050 7440 18106 7449
rect 17960 7404 18012 7410
rect 18050 7375 18106 7384
rect 17960 7346 18012 7352
rect 17972 6934 18000 7346
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17972 6458 18000 6870
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18156 6202 18184 8078
rect 18248 7313 18276 8298
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18340 7410 18368 8026
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18234 7304 18290 7313
rect 18432 7274 18460 17682
rect 18524 16250 18552 18022
rect 18616 17082 18644 18702
rect 18708 17338 18736 18838
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18616 17054 18736 17082
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 16590 18644 16934
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15570 18552 16050
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18616 12753 18644 16526
rect 18708 15094 18736 17054
rect 18800 16590 18828 18022
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18708 14600 18736 15030
rect 18788 14612 18840 14618
rect 18708 14572 18788 14600
rect 18788 14554 18840 14560
rect 18892 13977 18920 18634
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 18358 19472 18566
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19064 18216 19116 18222
rect 19168 18193 19196 18294
rect 19064 18158 19116 18164
rect 19154 18184 19210 18193
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18984 14074 19012 18090
rect 19076 17882 19104 18158
rect 19154 18119 19210 18128
rect 19430 18184 19486 18193
rect 19430 18119 19486 18128
rect 19444 18086 19472 18119
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19352 17762 19380 17818
rect 19076 17734 19380 17762
rect 19076 16182 19104 17734
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18878 13968 18934 13977
rect 18878 13903 18934 13912
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18234 7239 18290 7248
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18328 6928 18380 6934
rect 18328 6870 18380 6876
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6322 18276 6598
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18064 6174 18184 6202
rect 18236 6180 18288 6186
rect 18064 5574 18092 6174
rect 18236 6122 18288 6128
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18156 5098 18184 6054
rect 18248 5710 18276 6122
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18236 5160 18288 5166
rect 18236 5102 18288 5108
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17972 3534 18000 3878
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17880 3346 17908 3470
rect 17880 3318 18000 3346
rect 17972 3058 18000 3318
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17236 2650 17264 2926
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 1986 16436 2246
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16408 1958 16620 1986
rect 16592 800 16620 1958
rect 16960 800 16988 2314
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17328 800 17356 2246
rect 17696 800 17724 2246
rect 18064 800 18092 3606
rect 18156 3194 18184 4218
rect 18248 3670 18276 5102
rect 18236 3664 18288 3670
rect 18340 3641 18368 6870
rect 18432 6662 18460 6938
rect 18524 6730 18552 12038
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18616 11665 18644 11834
rect 18602 11656 18658 11665
rect 18602 11591 18658 11600
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18616 6934 18644 9415
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 8906 18828 8978
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18892 6798 18920 8774
rect 18984 8634 19012 14010
rect 19076 12986 19104 16118
rect 19536 15910 19564 21247
rect 20626 20904 20682 20913
rect 20626 20839 20682 20848
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19904 20262 19932 20402
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 20166 19816 20222 19825
rect 20166 19751 20222 19760
rect 20180 19718 20208 19751
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19628 17649 19656 18566
rect 19614 17640 19670 17649
rect 19614 17575 19670 17584
rect 19812 17270 19840 18702
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19904 16130 19932 17682
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19720 16102 19932 16130
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19536 14822 19564 15302
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 14414 19564 14758
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19352 14074 19380 14350
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19536 12986 19564 14350
rect 19720 14074 19748 16102
rect 19800 16040 19852 16046
rect 19892 16040 19944 16046
rect 19800 15982 19852 15988
rect 19890 16008 19892 16017
rect 19944 16008 19946 16017
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19076 11830 19104 12922
rect 19720 12918 19748 13874
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19812 12850 19840 15982
rect 19890 15943 19946 15952
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19628 11354 19656 12038
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19536 10062 19564 10542
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19430 9888 19486 9897
rect 19430 9823 19486 9832
rect 19444 9466 19472 9823
rect 19628 9654 19656 10746
rect 19720 10554 19748 12106
rect 19812 11778 19840 12786
rect 19904 12170 19932 15846
rect 19996 15042 20024 17478
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20088 16794 20116 17138
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19996 15014 20116 15042
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19996 12714 20024 14282
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19892 12164 19944 12170
rect 19892 12106 19944 12112
rect 19996 12102 20024 12650
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19812 11750 20024 11778
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19812 10742 19840 11562
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19720 10526 19840 10554
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19708 9512 19760 9518
rect 19444 9438 19656 9466
rect 19708 9454 19760 9460
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19628 9178 19656 9438
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19628 8974 19656 9114
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 19076 8022 19104 8502
rect 19720 8498 19748 9454
rect 19812 9110 19840 10526
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19904 9042 19932 11018
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18880 6792 18932 6798
rect 18786 6760 18842 6769
rect 18512 6724 18564 6730
rect 18880 6734 18932 6740
rect 18786 6695 18788 6704
rect 18512 6666 18564 6672
rect 18840 6695 18842 6704
rect 18788 6666 18840 6672
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18432 4049 18460 6598
rect 18510 6216 18566 6225
rect 18510 6151 18566 6160
rect 18524 5273 18552 6151
rect 18616 5914 18644 6598
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18418 4040 18474 4049
rect 18418 3975 18474 3984
rect 18236 3606 18288 3612
rect 18326 3632 18382 3641
rect 18326 3567 18382 3576
rect 18420 3596 18472 3602
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18340 2446 18368 3567
rect 18420 3538 18472 3544
rect 18432 2774 18460 3538
rect 18524 2961 18552 5199
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18616 4457 18644 5034
rect 18602 4448 18658 4457
rect 18602 4383 18658 4392
rect 18616 4282 18644 4383
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18708 4128 18736 6190
rect 18984 6186 19012 7414
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19076 7002 19104 7278
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 19536 6662 19564 7346
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19628 6322 19656 6598
rect 19720 6390 19748 8434
rect 19800 8356 19852 8362
rect 19800 8298 19852 8304
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18984 5386 19012 6122
rect 18616 4100 18736 4128
rect 18892 5358 19012 5386
rect 18616 3126 18644 4100
rect 18892 4078 18920 5358
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18708 3194 18736 3946
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18604 3120 18656 3126
rect 18656 3068 18736 3074
rect 18604 3062 18736 3068
rect 18616 3046 18736 3062
rect 18510 2952 18566 2961
rect 18510 2887 18566 2896
rect 18432 2746 18644 2774
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18432 800 18460 2518
rect 18616 2378 18644 2746
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18708 1737 18736 3046
rect 18694 1728 18750 1737
rect 18694 1663 18750 1672
rect 18800 800 18828 3946
rect 18892 3602 18920 4014
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18984 3505 19012 5170
rect 19076 5098 19104 6258
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19168 5166 19196 5510
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19720 4146 19748 5510
rect 19812 4622 19840 8298
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19338 4040 19394 4049
rect 19338 3975 19394 3984
rect 19352 3942 19380 3975
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18970 3496 19026 3505
rect 18892 3454 18970 3482
rect 18892 3058 18920 3454
rect 18970 3431 19026 3440
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18878 2952 18934 2961
rect 18878 2887 18934 2896
rect 18892 2446 18920 2887
rect 18984 2553 19012 3130
rect 18970 2544 19026 2553
rect 18970 2479 19026 2488
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 19076 1306 19104 3606
rect 19812 2990 19840 4558
rect 19904 4554 19932 8978
rect 19996 7886 20024 11750
rect 20088 10266 20116 15014
rect 20180 13410 20208 18770
rect 20272 16561 20300 20538
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 19281 20484 20198
rect 20640 20058 20668 20839
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20442 19272 20498 19281
rect 20442 19207 20498 19216
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18290 20392 18566
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17649 20484 18022
rect 20732 17678 20760 19790
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20720 17672 20772 17678
rect 20442 17640 20498 17649
rect 20720 17614 20772 17620
rect 20442 17575 20498 17584
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20258 16552 20314 16561
rect 20258 16487 20314 16496
rect 20364 16114 20392 16934
rect 20456 16658 20484 17478
rect 20640 16697 20668 17478
rect 20824 17338 20852 18838
rect 20916 18057 20944 19110
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 20996 18080 21048 18086
rect 20902 18048 20958 18057
rect 20996 18022 21048 18028
rect 20902 17983 20958 17992
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20626 16688 20682 16697
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20536 16652 20588 16658
rect 20626 16623 20682 16632
rect 20536 16594 20588 16600
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20364 14346 20392 15642
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20350 13560 20406 13569
rect 20350 13495 20406 13504
rect 20180 13382 20300 13410
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20180 12986 20208 13194
rect 20272 12986 20300 13382
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20180 11898 20208 12922
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20272 12322 20300 12786
rect 20364 12442 20392 13495
rect 20456 13297 20484 15302
rect 20442 13288 20498 13297
rect 20442 13223 20498 13232
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20272 12294 20392 12322
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20272 11830 20300 12174
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20258 11112 20314 11121
rect 20258 11047 20314 11056
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20088 9926 20116 10066
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 4706 20024 7686
rect 20088 7342 20116 9862
rect 20168 9104 20220 9110
rect 20168 9046 20220 9052
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20088 6322 20116 6802
rect 20180 6798 20208 9046
rect 20272 8974 20300 11047
rect 20364 10130 20392 12294
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8022 20300 8910
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20272 6610 20300 7822
rect 20364 7274 20392 9522
rect 20456 8090 20484 11698
rect 20548 11626 20576 16594
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 16182 20668 16526
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20732 15502 20760 16458
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20824 14822 20852 17070
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20640 14006 20668 14350
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20640 11150 20668 11834
rect 20732 11694 20760 14350
rect 20824 13258 20852 14758
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20640 10810 20668 11086
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20548 9110 20576 9590
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20548 7954 20576 8774
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20364 6866 20392 7210
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20180 6582 20300 6610
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 20088 4808 20116 6258
rect 20180 5574 20208 6582
rect 20364 6474 20392 6802
rect 20272 6446 20392 6474
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20272 5114 20300 6446
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20364 5914 20392 6258
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20272 5086 20392 5114
rect 20258 4992 20314 5001
rect 20258 4927 20314 4936
rect 20168 4820 20220 4826
rect 20088 4780 20168 4808
rect 20168 4762 20220 4768
rect 19996 4678 20208 4706
rect 19892 4548 19944 4554
rect 19892 4490 19944 4496
rect 19982 4176 20038 4185
rect 19982 4111 20038 4120
rect 19996 3058 20024 4111
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 20180 2446 20208 4678
rect 20272 4486 20300 4927
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 3534 20300 4422
rect 20364 4214 20392 5086
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20456 2650 20484 7686
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 7041 20576 7346
rect 20534 7032 20590 7041
rect 20534 6967 20590 6976
rect 20640 6662 20668 9862
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20732 6610 20760 11494
rect 20824 11082 20852 12242
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20824 10538 20852 11018
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20916 10146 20944 17478
rect 21008 15609 21036 18022
rect 21284 17882 21312 18226
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20994 15600 21050 15609
rect 20994 15535 21050 15544
rect 21100 15178 21128 16662
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21008 15150 21128 15178
rect 21008 13938 21036 15150
rect 21086 15056 21142 15065
rect 21086 14991 21142 15000
rect 21100 14618 21128 14991
rect 21192 14793 21220 16390
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21270 16008 21326 16017
rect 21270 15943 21272 15952
rect 21324 15943 21326 15952
rect 21272 15914 21324 15920
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21178 14784 21234 14793
rect 21178 14719 21234 14728
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21284 14414 21312 15302
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21272 14408 21324 14414
rect 21086 14376 21142 14385
rect 21272 14350 21324 14356
rect 21086 14311 21142 14320
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21100 13530 21128 14311
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 21008 12442 21036 12718
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11558 21036 12038
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 21284 11354 21312 12786
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 20916 10118 21036 10146
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20916 9722 20944 9862
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20824 6730 20852 8774
rect 21008 8090 21036 10118
rect 21284 9738 21312 11290
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21192 9710 21312 9738
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21192 7410 21220 9710
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 7546 21312 9522
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20904 6656 20956 6662
rect 20732 6604 20904 6610
rect 20732 6598 20956 6604
rect 20732 6582 20944 6598
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20548 5234 20576 5510
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20534 5128 20590 5137
rect 20534 5063 20536 5072
rect 20588 5063 20590 5072
rect 20536 5034 20588 5040
rect 20640 4146 20668 5850
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3194 20668 4082
rect 20732 3534 20760 5238
rect 20824 5166 20852 6582
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5302 20944 6054
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19076 1278 19196 1306
rect 19168 800 19196 1278
rect 19536 800 19564 2042
rect 19904 870 20024 898
rect 19904 800 19932 870
rect 15212 734 15424 762
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 19996 762 20024 870
rect 20180 762 20208 2382
rect 20260 2304 20312 2310
rect 20260 2246 20312 2252
rect 20272 800 20300 2246
rect 20640 800 20668 2994
rect 20824 2961 20852 5102
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4826 20944 4966
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20916 3602 20944 4762
rect 21008 4457 21036 6258
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5030 21128 6054
rect 21192 5846 21220 7346
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21376 6322 21404 6666
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 21192 4593 21220 5782
rect 21270 5264 21326 5273
rect 21270 5199 21326 5208
rect 21178 4584 21234 4593
rect 21178 4519 21234 4528
rect 20994 4448 21050 4457
rect 20994 4383 21050 4392
rect 21008 4185 21036 4383
rect 20994 4176 21050 4185
rect 20994 4111 21050 4120
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20810 2952 20866 2961
rect 20810 2887 20866 2896
rect 20916 2774 20944 3538
rect 21192 3534 21220 4519
rect 21284 4321 21312 5199
rect 21376 4486 21404 6258
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21270 4312 21326 4321
rect 21270 4247 21326 4256
rect 21284 4146 21312 4247
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21376 3777 21404 4422
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21376 3398 21404 3703
rect 21454 3496 21510 3505
rect 21454 3431 21510 3440
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21468 3194 21496 3431
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 20916 2746 21220 2774
rect 20994 2544 21050 2553
rect 21192 2514 21220 2746
rect 20994 2479 21050 2488
rect 21180 2508 21232 2514
rect 21008 2446 21036 2479
rect 21180 2450 21232 2456
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 21100 2009 21128 2246
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21086 2000 21142 2009
rect 21086 1935 21142 1944
rect 19996 734 20208 762
rect 20258 0 20314 800
rect 20626 0 20682 800
<< via2 >>
rect 3330 21256 3386 21312
rect 1950 20848 2006 20904
rect 2778 20440 2834 20496
rect 2870 20032 2926 20088
rect 1950 19660 1952 19680
rect 1952 19660 2004 19680
rect 2004 19660 2006 19680
rect 1950 19624 2006 19660
rect 1950 19236 2006 19272
rect 1950 19216 1952 19236
rect 1952 19216 2004 19236
rect 2004 19216 2006 19236
rect 1858 18808 1914 18864
rect 1490 17584 1546 17640
rect 1582 17176 1638 17232
rect 1950 17992 2006 18048
rect 1398 14728 1454 14784
rect 2134 16360 2190 16416
rect 2318 15580 2320 15600
rect 2320 15580 2372 15600
rect 2372 15580 2374 15600
rect 2318 15544 2374 15580
rect 2778 18400 2834 18456
rect 2778 16768 2834 16824
rect 1766 13504 1822 13560
rect 1950 13096 2006 13152
rect 1582 8200 1638 8256
rect 1582 7812 1638 7848
rect 1582 7792 1584 7812
rect 1584 7792 1636 7812
rect 1636 7792 1638 7812
rect 1398 3712 1454 3768
rect 1766 3304 1822 3360
rect 2318 11736 2374 11792
rect 2134 5344 2190 5400
rect 1950 4936 2006 4992
rect 2134 3984 2190 4040
rect 1858 2080 1914 2136
rect 2962 16496 3018 16552
rect 2870 15952 2926 16008
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 2962 15136 3018 15192
rect 2778 14320 2834 14376
rect 2870 12144 2926 12200
rect 3054 12416 3110 12472
rect 3330 13912 3386 13968
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3146 11872 3202 11928
rect 3054 11464 3110 11520
rect 2594 5480 2650 5536
rect 2778 4528 2834 4584
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 4158 16652 4214 16688
rect 4158 16632 4160 16652
rect 4160 16632 4212 16652
rect 4212 16632 4214 16652
rect 4066 12688 4122 12744
rect 4434 13232 4490 13288
rect 4066 12300 4122 12336
rect 4066 12280 4068 12300
rect 4068 12280 4120 12300
rect 4120 12280 4122 12300
rect 3882 10104 3938 10160
rect 3330 9152 3386 9208
rect 3146 6568 3202 6624
rect 3054 5344 3110 5400
rect 2870 4120 2926 4176
rect 3606 9560 3662 9616
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 4342 11076 4398 11112
rect 4342 11056 4344 11076
rect 4344 11056 4396 11076
rect 4396 11056 4398 11076
rect 4066 10512 4122 10568
rect 4066 9832 4122 9888
rect 4158 9424 4214 9480
rect 4066 8608 4122 8664
rect 4250 8336 4306 8392
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3330 2896 3386 2952
rect 3238 2488 3294 2544
rect 3790 6160 3846 6216
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3974 7520 4030 7576
rect 4526 6840 4582 6896
rect 4066 6432 4122 6488
rect 3974 6296 4030 6352
rect 3974 6196 3976 6216
rect 3976 6196 4028 6216
rect 4028 6196 4030 6216
rect 3974 6160 4030 6196
rect 4066 4684 4122 4720
rect 4066 4664 4068 4684
rect 4068 4664 4120 4684
rect 4120 4664 4122 4684
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 7102 19352 7158 19408
rect 5538 18264 5594 18320
rect 5354 17076 5356 17096
rect 5356 17076 5408 17096
rect 5408 17076 5410 17096
rect 5354 17040 5410 17076
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 5722 17992 5778 18048
rect 5170 14728 5226 14784
rect 4894 10648 4950 10704
rect 4710 9424 4766 9480
rect 4434 4564 4436 4584
rect 4436 4564 4488 4584
rect 4488 4564 4490 4584
rect 4434 4528 4490 4564
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 1672 3478 1728
rect 4894 7828 4896 7848
rect 4896 7828 4948 7848
rect 4948 7828 4950 7848
rect 4894 7792 4950 7828
rect 5630 14456 5686 14512
rect 5630 12552 5686 12608
rect 5446 7384 5502 7440
rect 5170 4120 5226 4176
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5998 16632 6054 16688
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6550 15816 6606 15872
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5998 12724 6000 12744
rect 6000 12724 6052 12744
rect 6052 12724 6054 12744
rect 5998 12688 6054 12724
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 7470 17584 7526 17640
rect 6918 15952 6974 16008
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6090 9968 6146 10024
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5722 5616 5778 5672
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6918 11056 6974 11112
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6458 5616 6514 5672
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 7102 12044 7104 12064
rect 7104 12044 7156 12064
rect 7156 12044 7158 12064
rect 7102 12008 7158 12044
rect 7746 16496 7802 16552
rect 7562 13368 7618 13424
rect 6826 7248 6882 7304
rect 6642 5344 6698 5400
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5538 3596 5594 3632
rect 5538 3576 5540 3596
rect 5540 3576 5592 3596
rect 5592 3576 5594 3596
rect 5814 3032 5870 3088
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6734 3168 6790 3224
rect 7010 3304 7066 3360
rect 6918 2488 6974 2544
rect 8022 16632 8078 16688
rect 7746 10784 7802 10840
rect 7654 8084 7710 8120
rect 7654 8064 7656 8084
rect 7656 8064 7708 8084
rect 7708 8064 7710 8084
rect 7930 10784 7986 10840
rect 7930 9968 7986 10024
rect 8206 14728 8262 14784
rect 8206 12044 8208 12064
rect 8208 12044 8260 12064
rect 8260 12044 8262 12064
rect 8206 12008 8262 12044
rect 8206 8880 8262 8936
rect 8022 5480 8078 5536
rect 7746 2896 7802 2952
rect 7930 3984 7986 4040
rect 9954 19352 10010 19408
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9034 9424 9090 9480
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9310 7248 9366 7304
rect 8850 6332 8852 6352
rect 8852 6332 8904 6352
rect 8904 6332 8906 6352
rect 8850 6296 8906 6332
rect 8758 6160 8814 6216
rect 8942 6180 8998 6216
rect 8942 6160 8944 6180
rect 8944 6160 8996 6180
rect 8996 6160 8998 6180
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9678 12824 9734 12880
rect 10138 17992 10194 18048
rect 9678 12280 9734 12336
rect 9586 6840 9642 6896
rect 9586 6296 9642 6352
rect 10138 11756 10194 11792
rect 10138 11736 10140 11756
rect 10140 11736 10192 11756
rect 10192 11736 10194 11756
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 11058 19660 11060 19680
rect 11060 19660 11112 19680
rect 11112 19660 11114 19680
rect 11058 19624 11114 19660
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11610 18808 11666 18864
rect 10506 13232 10562 13288
rect 10414 12688 10470 12744
rect 9862 7928 9918 7984
rect 9310 5616 9366 5672
rect 9678 5616 9734 5672
rect 8942 4140 8998 4176
rect 8942 4120 8944 4140
rect 8944 4120 8996 4140
rect 8996 4120 8998 4140
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9402 4120 9458 4176
rect 9310 4004 9366 4040
rect 9310 3984 9312 4004
rect 9312 3984 9364 4004
rect 9364 3984 9366 4004
rect 9586 4020 9588 4040
rect 9588 4020 9640 4040
rect 9640 4020 9642 4040
rect 9586 3984 9642 4020
rect 8942 3440 8998 3496
rect 9218 3304 9274 3360
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9770 2796 9772 2816
rect 9772 2796 9824 2816
rect 9824 2796 9826 2816
rect 9770 2760 9826 2796
rect 11058 18264 11114 18320
rect 10966 16652 11022 16688
rect 10966 16632 10968 16652
rect 10968 16632 11020 16652
rect 11020 16632 11022 16652
rect 10782 16088 10838 16144
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 12622 18672 12678 18728
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10690 10512 10746 10568
rect 10598 9968 10654 10024
rect 10322 8200 10378 8256
rect 10322 7792 10378 7848
rect 10230 2760 10286 2816
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10966 7248 11022 7304
rect 11058 5344 11114 5400
rect 10782 4664 10838 4720
rect 10690 3848 10746 3904
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11150 3848 11206 3904
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11334 3884 11336 3904
rect 11336 3884 11388 3904
rect 11388 3884 11390 3904
rect 11334 3848 11390 3884
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12162 10104 12218 10160
rect 12254 8880 12310 8936
rect 13174 12688 13230 12744
rect 13542 15408 13598 15464
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13082 8200 13138 8256
rect 13082 4140 13138 4176
rect 13082 4120 13084 4140
rect 13084 4120 13136 4140
rect 13136 4120 13138 4140
rect 13266 3576 13322 3632
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14278 11600 14334 11656
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13818 3712 13874 3768
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 14646 11056 14702 11112
rect 14462 3032 14518 3088
rect 16946 18808 17002 18864
rect 19522 21256 19578 21312
rect 18050 20440 18106 20496
rect 17958 19932 17960 19952
rect 17960 19932 18012 19952
rect 18012 19932 18014 19952
rect 17958 19896 18014 19932
rect 17498 19352 17554 19408
rect 15290 16632 15346 16688
rect 15382 15000 15438 15056
rect 17406 18808 17462 18864
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16486 18128 16542 18184
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 13818 2896 13874 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15382 4256 15438 4312
rect 15934 6332 15936 6352
rect 15936 6332 15988 6352
rect 15988 6332 15990 6352
rect 15934 6296 15990 6332
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16578 5228 16634 5264
rect 16578 5208 16580 5228
rect 16580 5208 16632 5228
rect 16632 5208 16634 5228
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16670 3612 16672 3632
rect 16672 3612 16724 3632
rect 16724 3612 16726 3632
rect 16670 3576 16726 3612
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17038 6160 17094 6216
rect 17774 18264 17830 18320
rect 17498 7384 17554 7440
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 18050 17212 18052 17232
rect 18052 17212 18104 17232
rect 18104 17212 18106 17232
rect 18050 17176 18106 17212
rect 17958 16632 18014 16688
rect 18234 18708 18236 18728
rect 18236 18708 18288 18728
rect 18288 18708 18290 18728
rect 18234 18672 18290 18708
rect 18234 16088 18290 16144
rect 18050 12280 18106 12336
rect 18050 11756 18106 11792
rect 18050 11736 18052 11756
rect 18052 11736 18104 11756
rect 18104 11736 18106 11756
rect 17958 9968 18014 10024
rect 17958 9016 18014 9072
rect 18142 8472 18198 8528
rect 17774 7792 17830 7848
rect 17682 6568 17738 6624
rect 17314 5616 17370 5672
rect 17774 4120 17830 4176
rect 18050 7384 18106 7440
rect 18234 7248 18290 7304
rect 19154 18128 19210 18184
rect 19430 18128 19486 18184
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 18878 13912 18934 13968
rect 18602 12688 18658 12744
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 18602 11600 18658 11656
rect 18602 9424 18658 9480
rect 20626 20848 20682 20904
rect 20166 19760 20222 19816
rect 19614 17584 19670 17640
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19890 15988 19892 16008
rect 19892 15988 19944 16008
rect 19944 15988 19946 16008
rect 19890 15952 19946 15988
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19430 9832 19486 9888
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 18786 6724 18842 6760
rect 18786 6704 18788 6724
rect 18788 6704 18840 6724
rect 18840 6704 18842 6724
rect 18510 6160 18566 6216
rect 18510 5208 18566 5264
rect 18418 3984 18474 4040
rect 18326 3576 18382 3632
rect 18602 4392 18658 4448
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18510 2896 18566 2952
rect 18694 1672 18750 1728
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19338 3984 19394 4040
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 18970 3440 19026 3496
rect 18878 2896 18934 2952
rect 18970 2488 19026 2544
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 20442 19216 20498 19272
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 20442 17584 20498 17640
rect 20258 16496 20314 16552
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 20902 17992 20958 18048
rect 20626 16632 20682 16688
rect 20350 13504 20406 13560
rect 20442 13232 20498 13288
rect 20258 11056 20314 11112
rect 20258 4936 20314 4992
rect 19982 4120 20038 4176
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20534 6976 20590 7032
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 20994 15544 21050 15600
rect 21086 15000 21142 15056
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21270 15972 21326 16008
rect 21270 15952 21272 15972
rect 21272 15952 21324 15972
rect 21324 15952 21326 15972
rect 21178 14728 21234 14784
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21086 14320 21142 14376
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 20534 5092 20590 5128
rect 20534 5072 20536 5092
rect 20536 5072 20588 5092
rect 20588 5072 20590 5092
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21270 5208 21326 5264
rect 21178 4528 21234 4584
rect 20994 4392 21050 4448
rect 20994 4120 21050 4176
rect 20810 2896 20866 2952
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21270 4256 21326 4312
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21362 3712 21418 3768
rect 21454 3440 21510 3496
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 20994 2488 21050 2544
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21086 1944 21142 2000
<< metal3 >>
rect 0 21314 800 21344
rect 3325 21314 3391 21317
rect 0 21312 3391 21314
rect 0 21256 3330 21312
rect 3386 21256 3391 21312
rect 0 21254 3391 21256
rect 0 21224 800 21254
rect 3325 21251 3391 21254
rect 19517 21314 19583 21317
rect 22200 21314 23000 21344
rect 19517 21312 23000 21314
rect 19517 21256 19522 21312
rect 19578 21256 23000 21312
rect 19517 21254 23000 21256
rect 19517 21251 19583 21254
rect 22200 21224 23000 21254
rect 0 20906 800 20936
rect 1945 20906 2011 20909
rect 0 20904 2011 20906
rect 0 20848 1950 20904
rect 2006 20848 2011 20904
rect 0 20846 2011 20848
rect 0 20816 800 20846
rect 1945 20843 2011 20846
rect 20621 20906 20687 20909
rect 22200 20906 23000 20936
rect 20621 20904 23000 20906
rect 20621 20848 20626 20904
rect 20682 20848 23000 20904
rect 20621 20846 23000 20848
rect 20621 20843 20687 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 2773 20498 2839 20501
rect 0 20496 2839 20498
rect 0 20440 2778 20496
rect 2834 20440 2839 20496
rect 0 20438 2839 20440
rect 0 20408 800 20438
rect 2773 20435 2839 20438
rect 18045 20498 18111 20501
rect 22200 20498 23000 20528
rect 18045 20496 23000 20498
rect 18045 20440 18050 20496
rect 18106 20440 23000 20496
rect 18045 20438 23000 20440
rect 18045 20435 18111 20438
rect 22200 20408 23000 20438
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 2865 20090 2931 20093
rect 22200 20090 23000 20120
rect 0 20088 2931 20090
rect 0 20032 2870 20088
rect 2926 20032 2931 20088
rect 0 20030 2931 20032
rect 0 20000 800 20030
rect 2865 20027 2931 20030
rect 19566 20030 23000 20090
rect 17953 19954 18019 19957
rect 19566 19954 19626 20030
rect 22200 20000 23000 20030
rect 17953 19952 19626 19954
rect 17953 19896 17958 19952
rect 18014 19896 19626 19952
rect 17953 19894 19626 19896
rect 17953 19891 18019 19894
rect 20161 19818 20227 19821
rect 20161 19816 22202 19818
rect 20161 19760 20166 19816
rect 20222 19760 22202 19816
rect 20161 19758 22202 19760
rect 20161 19755 20227 19758
rect 22142 19712 22202 19758
rect 0 19682 800 19712
rect 1945 19682 2011 19685
rect 11053 19684 11119 19685
rect 11053 19682 11100 19684
rect 0 19680 2011 19682
rect 0 19624 1950 19680
rect 2006 19624 2011 19680
rect 0 19622 2011 19624
rect 11008 19680 11100 19682
rect 11008 19624 11058 19680
rect 11008 19622 11100 19624
rect 0 19592 800 19622
rect 1945 19619 2011 19622
rect 11053 19620 11100 19622
rect 11164 19620 11170 19684
rect 22142 19622 23000 19712
rect 11053 19619 11119 19620
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 3366 19348 3372 19412
rect 3436 19410 3442 19412
rect 7097 19410 7163 19413
rect 3436 19408 7163 19410
rect 3436 19352 7102 19408
rect 7158 19352 7163 19408
rect 3436 19350 7163 19352
rect 3436 19348 3442 19350
rect 7097 19347 7163 19350
rect 9254 19348 9260 19412
rect 9324 19410 9330 19412
rect 9949 19410 10015 19413
rect 9324 19408 10015 19410
rect 9324 19352 9954 19408
rect 10010 19352 10015 19408
rect 9324 19350 10015 19352
rect 9324 19348 9330 19350
rect 9949 19347 10015 19350
rect 16982 19348 16988 19412
rect 17052 19410 17058 19412
rect 17493 19410 17559 19413
rect 17052 19408 17559 19410
rect 17052 19352 17498 19408
rect 17554 19352 17559 19408
rect 17052 19350 17559 19352
rect 17052 19348 17058 19350
rect 17493 19347 17559 19350
rect 0 19274 800 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 800 19214
rect 1945 19211 2011 19214
rect 20437 19274 20503 19277
rect 22200 19274 23000 19304
rect 20437 19272 23000 19274
rect 20437 19216 20442 19272
rect 20498 19216 23000 19272
rect 20437 19214 23000 19216
rect 20437 19211 20503 19214
rect 22200 19184 23000 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 1853 18866 1919 18869
rect 0 18864 1919 18866
rect 0 18808 1858 18864
rect 1914 18808 1919 18864
rect 0 18806 1919 18808
rect 0 18776 800 18806
rect 1853 18803 1919 18806
rect 11605 18866 11671 18869
rect 16941 18866 17007 18869
rect 11605 18864 17007 18866
rect 11605 18808 11610 18864
rect 11666 18808 16946 18864
rect 17002 18808 17007 18864
rect 11605 18806 17007 18808
rect 11605 18803 11671 18806
rect 16941 18803 17007 18806
rect 17401 18866 17467 18869
rect 22200 18866 23000 18896
rect 17401 18864 23000 18866
rect 17401 18808 17406 18864
rect 17462 18808 23000 18864
rect 17401 18806 23000 18808
rect 17401 18803 17467 18806
rect 22200 18776 23000 18806
rect 12617 18730 12683 18733
rect 18229 18730 18295 18733
rect 12617 18728 18295 18730
rect 12617 18672 12622 18728
rect 12678 18672 18234 18728
rect 18290 18672 18295 18728
rect 12617 18670 18295 18672
rect 12617 18667 12683 18670
rect 18229 18667 18295 18670
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 2773 18458 2839 18461
rect 22200 18458 23000 18488
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18368 800 18398
rect 2773 18395 2839 18398
rect 22142 18368 23000 18458
rect 5533 18322 5599 18325
rect 11053 18322 11119 18325
rect 5533 18320 11119 18322
rect 5533 18264 5538 18320
rect 5594 18264 11058 18320
rect 11114 18264 11119 18320
rect 5533 18262 11119 18264
rect 5533 18259 5599 18262
rect 11053 18259 11119 18262
rect 17769 18322 17835 18325
rect 22142 18322 22202 18368
rect 17769 18320 22202 18322
rect 17769 18264 17774 18320
rect 17830 18264 22202 18320
rect 17769 18262 22202 18264
rect 17769 18259 17835 18262
rect 16481 18186 16547 18189
rect 19149 18186 19215 18189
rect 16481 18184 19215 18186
rect 16481 18128 16486 18184
rect 16542 18128 19154 18184
rect 19210 18128 19215 18184
rect 16481 18126 19215 18128
rect 16481 18123 16547 18126
rect 19149 18123 19215 18126
rect 19425 18186 19491 18189
rect 19558 18186 19564 18188
rect 19425 18184 19564 18186
rect 19425 18128 19430 18184
rect 19486 18128 19564 18184
rect 19425 18126 19564 18128
rect 19425 18123 19491 18126
rect 19558 18124 19564 18126
rect 19628 18124 19634 18188
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 5206 17988 5212 18052
rect 5276 18050 5282 18052
rect 5717 18050 5783 18053
rect 10133 18052 10199 18053
rect 10133 18050 10180 18052
rect 5276 18048 5783 18050
rect 5276 17992 5722 18048
rect 5778 17992 5783 18048
rect 5276 17990 5783 17992
rect 10088 18048 10180 18050
rect 10088 17992 10138 18048
rect 10088 17990 10180 17992
rect 5276 17988 5282 17990
rect 5717 17987 5783 17990
rect 10133 17988 10180 17990
rect 10244 17988 10250 18052
rect 20897 18050 20963 18053
rect 22200 18050 23000 18080
rect 20897 18048 23000 18050
rect 20897 17992 20902 18048
rect 20958 17992 23000 18048
rect 20897 17990 23000 17992
rect 10133 17987 10199 17988
rect 20897 17987 20963 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 0 17642 800 17672
rect 1485 17642 1551 17645
rect 0 17640 1551 17642
rect 0 17584 1490 17640
rect 1546 17584 1551 17640
rect 0 17582 1551 17584
rect 0 17552 800 17582
rect 1485 17579 1551 17582
rect 7465 17642 7531 17645
rect 19609 17642 19675 17645
rect 7465 17640 19675 17642
rect 7465 17584 7470 17640
rect 7526 17584 19614 17640
rect 19670 17584 19675 17640
rect 7465 17582 19675 17584
rect 7465 17579 7531 17582
rect 19609 17579 19675 17582
rect 20437 17642 20503 17645
rect 22200 17642 23000 17672
rect 20437 17640 23000 17642
rect 20437 17584 20442 17640
rect 20498 17584 23000 17640
rect 20437 17582 23000 17584
rect 20437 17579 20503 17582
rect 22200 17552 23000 17582
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1577 17234 1643 17237
rect 0 17232 1643 17234
rect 0 17176 1582 17232
rect 1638 17176 1643 17232
rect 0 17174 1643 17176
rect 0 17144 800 17174
rect 1577 17171 1643 17174
rect 18045 17234 18111 17237
rect 22200 17234 23000 17264
rect 18045 17232 23000 17234
rect 18045 17176 18050 17232
rect 18106 17176 23000 17232
rect 18045 17174 23000 17176
rect 18045 17171 18111 17174
rect 22200 17144 23000 17174
rect 5349 17098 5415 17101
rect 10542 17098 10548 17100
rect 5349 17096 10548 17098
rect 5349 17040 5354 17096
rect 5410 17040 10548 17096
rect 5349 17038 10548 17040
rect 5349 17035 5415 17038
rect 10542 17036 10548 17038
rect 10612 17036 10618 17100
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 2773 16826 2839 16829
rect 22200 16826 23000 16856
rect 0 16824 2839 16826
rect 0 16768 2778 16824
rect 2834 16768 2839 16824
rect 0 16766 2839 16768
rect 0 16736 800 16766
rect 2773 16763 2839 16766
rect 19566 16766 23000 16826
rect 4153 16690 4219 16693
rect 4286 16690 4292 16692
rect 4153 16688 4292 16690
rect 4153 16632 4158 16688
rect 4214 16632 4292 16688
rect 4153 16630 4292 16632
rect 4153 16627 4219 16630
rect 4286 16628 4292 16630
rect 4356 16628 4362 16692
rect 5993 16690 6059 16693
rect 6678 16690 6684 16692
rect 5993 16688 6684 16690
rect 5993 16632 5998 16688
rect 6054 16632 6684 16688
rect 5993 16630 6684 16632
rect 5993 16627 6059 16630
rect 6678 16628 6684 16630
rect 6748 16628 6754 16692
rect 8017 16690 8083 16693
rect 8150 16690 8156 16692
rect 8017 16688 8156 16690
rect 8017 16632 8022 16688
rect 8078 16632 8156 16688
rect 8017 16630 8156 16632
rect 8017 16627 8083 16630
rect 8150 16628 8156 16630
rect 8220 16628 8226 16692
rect 10961 16690 11027 16693
rect 15285 16690 15351 16693
rect 10961 16688 15351 16690
rect 10961 16632 10966 16688
rect 11022 16632 15290 16688
rect 15346 16632 15351 16688
rect 10961 16630 15351 16632
rect 10961 16627 11027 16630
rect 15285 16627 15351 16630
rect 17953 16690 18019 16693
rect 19566 16690 19626 16766
rect 22200 16736 23000 16766
rect 17953 16688 19626 16690
rect 17953 16632 17958 16688
rect 18014 16632 19626 16688
rect 17953 16630 19626 16632
rect 17953 16627 18019 16630
rect 20478 16628 20484 16692
rect 20548 16690 20554 16692
rect 20621 16690 20687 16693
rect 20548 16688 20687 16690
rect 20548 16632 20626 16688
rect 20682 16632 20687 16688
rect 20548 16630 20687 16632
rect 20548 16628 20554 16630
rect 20621 16627 20687 16630
rect 2957 16554 3023 16557
rect 7741 16554 7807 16557
rect 2957 16552 7807 16554
rect 2957 16496 2962 16552
rect 3018 16496 7746 16552
rect 7802 16496 7807 16552
rect 2957 16494 7807 16496
rect 2957 16491 3023 16494
rect 7741 16491 7807 16494
rect 20253 16554 20319 16557
rect 20253 16552 22202 16554
rect 20253 16496 20258 16552
rect 20314 16496 22202 16552
rect 20253 16494 22202 16496
rect 20253 16491 20319 16494
rect 22142 16448 22202 16494
rect 0 16418 800 16448
rect 2129 16418 2195 16421
rect 0 16416 2195 16418
rect 0 16360 2134 16416
rect 2190 16360 2195 16416
rect 0 16358 2195 16360
rect 22142 16358 23000 16448
rect 0 16328 800 16358
rect 2129 16355 2195 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 10777 16146 10843 16149
rect 18229 16146 18295 16149
rect 10777 16144 18295 16146
rect 10777 16088 10782 16144
rect 10838 16088 18234 16144
rect 18290 16088 18295 16144
rect 10777 16086 18295 16088
rect 10777 16083 10843 16086
rect 18229 16083 18295 16086
rect 0 16010 800 16040
rect 2865 16010 2931 16013
rect 0 16008 2931 16010
rect 0 15952 2870 16008
rect 2926 15952 2931 16008
rect 0 15950 2931 15952
rect 0 15920 800 15950
rect 2865 15947 2931 15950
rect 6913 16010 6979 16013
rect 7046 16010 7052 16012
rect 6913 16008 7052 16010
rect 6913 15952 6918 16008
rect 6974 15952 7052 16008
rect 6913 15950 7052 15952
rect 6913 15947 6979 15950
rect 7046 15948 7052 15950
rect 7116 15948 7122 16012
rect 19885 16010 19951 16013
rect 7238 16008 19951 16010
rect 7238 15952 19890 16008
rect 19946 15952 19951 16008
rect 7238 15950 19951 15952
rect 6545 15874 6611 15877
rect 7238 15874 7298 15950
rect 19885 15947 19951 15950
rect 21265 16010 21331 16013
rect 22200 16010 23000 16040
rect 21265 16008 23000 16010
rect 21265 15952 21270 16008
rect 21326 15952 23000 16008
rect 21265 15950 23000 15952
rect 21265 15947 21331 15950
rect 22200 15920 23000 15950
rect 6545 15872 7298 15874
rect 6545 15816 6550 15872
rect 6606 15816 7298 15872
rect 6545 15814 7298 15816
rect 6545 15811 6611 15814
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 2313 15602 2379 15605
rect 0 15600 2379 15602
rect 0 15544 2318 15600
rect 2374 15544 2379 15600
rect 0 15542 2379 15544
rect 0 15512 800 15542
rect 2313 15539 2379 15542
rect 20989 15602 21055 15605
rect 22200 15602 23000 15632
rect 20989 15600 23000 15602
rect 20989 15544 20994 15600
rect 21050 15544 23000 15600
rect 20989 15542 23000 15544
rect 20989 15539 21055 15542
rect 22200 15512 23000 15542
rect 9438 15404 9444 15468
rect 9508 15466 9514 15468
rect 13537 15466 13603 15469
rect 9508 15464 13603 15466
rect 9508 15408 13542 15464
rect 13598 15408 13603 15464
rect 9508 15406 13603 15408
rect 9508 15404 9514 15406
rect 13537 15403 13603 15406
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 2957 15194 3023 15197
rect 22200 15194 23000 15224
rect 0 15192 3023 15194
rect 0 15136 2962 15192
rect 3018 15136 3023 15192
rect 0 15134 3023 15136
rect 0 15104 800 15134
rect 2957 15131 3023 15134
rect 22142 15104 23000 15194
rect 15377 15058 15443 15061
rect 16982 15058 16988 15060
rect 15377 15056 16988 15058
rect 15377 15000 15382 15056
rect 15438 15000 16988 15056
rect 15377 14998 16988 15000
rect 15377 14995 15443 14998
rect 16982 14996 16988 14998
rect 17052 14996 17058 15060
rect 21081 15058 21147 15061
rect 22142 15058 22202 15104
rect 21081 15056 22202 15058
rect 21081 15000 21086 15056
rect 21142 15000 22202 15056
rect 21081 14998 22202 15000
rect 21081 14995 21147 14998
rect 0 14786 800 14816
rect 1393 14786 1459 14789
rect 0 14784 1459 14786
rect 0 14728 1398 14784
rect 1454 14728 1459 14784
rect 0 14726 1459 14728
rect 0 14696 800 14726
rect 1393 14723 1459 14726
rect 5165 14786 5231 14789
rect 8201 14786 8267 14789
rect 5165 14784 8267 14786
rect 5165 14728 5170 14784
rect 5226 14728 8206 14784
rect 8262 14728 8267 14784
rect 5165 14726 8267 14728
rect 5165 14723 5231 14726
rect 8201 14723 8267 14726
rect 21173 14786 21239 14789
rect 22200 14786 23000 14816
rect 21173 14784 23000 14786
rect 21173 14728 21178 14784
rect 21234 14728 23000 14784
rect 21173 14726 23000 14728
rect 21173 14723 21239 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 5625 14514 5691 14517
rect 5582 14512 5691 14514
rect 5582 14456 5630 14512
rect 5686 14456 5691 14512
rect 5582 14451 5691 14456
rect 0 14378 800 14408
rect 2773 14378 2839 14381
rect 0 14376 2839 14378
rect 0 14320 2778 14376
rect 2834 14320 2839 14376
rect 0 14318 2839 14320
rect 0 14288 800 14318
rect 2773 14315 2839 14318
rect 0 13970 800 14000
rect 3325 13970 3391 13973
rect 0 13968 3391 13970
rect 0 13912 3330 13968
rect 3386 13912 3391 13968
rect 0 13910 3391 13912
rect 0 13880 800 13910
rect 3325 13907 3391 13910
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 1761 13562 1827 13565
rect 0 13560 1827 13562
rect 0 13504 1766 13560
rect 1822 13504 1827 13560
rect 0 13502 1827 13504
rect 0 13472 800 13502
rect 1761 13499 1827 13502
rect 2814 13364 2820 13428
rect 2884 13426 2890 13428
rect 5582 13426 5642 14451
rect 21081 14378 21147 14381
rect 22200 14378 23000 14408
rect 21081 14376 23000 14378
rect 21081 14320 21086 14376
rect 21142 14320 23000 14376
rect 21081 14318 23000 14320
rect 21081 14315 21147 14318
rect 22200 14288 23000 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 18873 13970 18939 13973
rect 22200 13970 23000 14000
rect 18873 13968 23000 13970
rect 18873 13912 18878 13968
rect 18934 13912 23000 13968
rect 18873 13910 23000 13912
rect 18873 13907 18939 13910
rect 22200 13880 23000 13910
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 20345 13562 20411 13565
rect 22200 13562 23000 13592
rect 20345 13560 23000 13562
rect 20345 13504 20350 13560
rect 20406 13504 23000 13560
rect 20345 13502 23000 13504
rect 20345 13499 20411 13502
rect 22200 13472 23000 13502
rect 2884 13366 5642 13426
rect 7557 13426 7623 13429
rect 9622 13426 9628 13428
rect 7557 13424 9628 13426
rect 7557 13368 7562 13424
rect 7618 13368 9628 13424
rect 7557 13366 9628 13368
rect 2884 13364 2890 13366
rect 7557 13363 7623 13366
rect 9622 13364 9628 13366
rect 9692 13364 9698 13428
rect 4429 13290 4495 13293
rect 10501 13290 10567 13293
rect 4429 13288 10567 13290
rect 4429 13232 4434 13288
rect 4490 13232 10506 13288
rect 10562 13232 10567 13288
rect 4429 13230 10567 13232
rect 4429 13227 4495 13230
rect 10501 13227 10567 13230
rect 20437 13290 20503 13293
rect 20437 13288 22202 13290
rect 20437 13232 20442 13288
rect 20498 13232 22202 13288
rect 20437 13230 22202 13232
rect 20437 13227 20503 13230
rect 22142 13184 22202 13230
rect 0 13154 800 13184
rect 1945 13154 2011 13157
rect 0 13152 2011 13154
rect 0 13096 1950 13152
rect 2006 13096 2011 13152
rect 0 13094 2011 13096
rect 22142 13094 23000 13184
rect 0 13064 800 13094
rect 1945 13091 2011 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 8334 12820 8340 12884
rect 8404 12882 8410 12884
rect 9673 12882 9739 12885
rect 8404 12880 9739 12882
rect 8404 12824 9678 12880
rect 9734 12824 9739 12880
rect 8404 12822 9739 12824
rect 8404 12820 8410 12822
rect 9673 12819 9739 12822
rect 0 12746 800 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 800 12686
rect 4061 12683 4127 12686
rect 5993 12746 6059 12749
rect 10409 12746 10475 12749
rect 5993 12744 10475 12746
rect 5993 12688 5998 12744
rect 6054 12688 10414 12744
rect 10470 12688 10475 12744
rect 5993 12686 10475 12688
rect 5993 12683 6059 12686
rect 10409 12683 10475 12686
rect 10542 12684 10548 12748
rect 10612 12746 10618 12748
rect 13169 12746 13235 12749
rect 10612 12744 13235 12746
rect 10612 12688 13174 12744
rect 13230 12688 13235 12744
rect 10612 12686 13235 12688
rect 10612 12684 10618 12686
rect 13169 12683 13235 12686
rect 18597 12746 18663 12749
rect 22200 12746 23000 12776
rect 18597 12744 23000 12746
rect 18597 12688 18602 12744
rect 18658 12688 23000 12744
rect 18597 12686 23000 12688
rect 18597 12683 18663 12686
rect 22200 12656 23000 12686
rect 5625 12610 5691 12613
rect 5758 12610 5764 12612
rect 5625 12608 5764 12610
rect 5625 12552 5630 12608
rect 5686 12552 5764 12608
rect 5625 12550 5764 12552
rect 5625 12547 5691 12550
rect 5758 12548 5764 12550
rect 5828 12548 5834 12612
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 3049 12474 3115 12477
rect 3006 12472 3115 12474
rect 3006 12416 3054 12472
rect 3110 12416 3115 12472
rect 3006 12411 3115 12416
rect 0 12338 800 12368
rect 3006 12338 3066 12411
rect 0 12278 3066 12338
rect 4061 12338 4127 12341
rect 4286 12338 4292 12340
rect 4061 12336 4292 12338
rect 4061 12280 4066 12336
rect 4122 12280 4292 12336
rect 4061 12278 4292 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 4286 12276 4292 12278
rect 4356 12276 4362 12340
rect 4470 12276 4476 12340
rect 4540 12338 4546 12340
rect 8334 12338 8340 12340
rect 4540 12278 8340 12338
rect 4540 12276 4546 12278
rect 8334 12276 8340 12278
rect 8404 12276 8410 12340
rect 9673 12338 9739 12341
rect 9806 12338 9812 12340
rect 9673 12336 9812 12338
rect 9673 12280 9678 12336
rect 9734 12280 9812 12336
rect 9673 12278 9812 12280
rect 9673 12275 9739 12278
rect 9806 12276 9812 12278
rect 9876 12276 9882 12340
rect 18045 12338 18111 12341
rect 22200 12338 23000 12368
rect 18045 12336 23000 12338
rect 18045 12280 18050 12336
rect 18106 12280 23000 12336
rect 18045 12278 23000 12280
rect 18045 12275 18111 12278
rect 22200 12248 23000 12278
rect 2865 12202 2931 12205
rect 2865 12200 6746 12202
rect 2865 12144 2870 12200
rect 2926 12144 6746 12200
rect 2865 12142 6746 12144
rect 2865 12139 2931 12142
rect 6686 12066 6746 12142
rect 7097 12066 7163 12069
rect 7230 12066 7236 12068
rect 6686 12064 7236 12066
rect 6686 12008 7102 12064
rect 7158 12008 7236 12064
rect 6686 12006 7236 12008
rect 7097 12003 7163 12006
rect 7230 12004 7236 12006
rect 7300 12066 7306 12068
rect 8201 12066 8267 12069
rect 7300 12064 8267 12066
rect 7300 12008 8206 12064
rect 8262 12008 8267 12064
rect 7300 12006 8267 12008
rect 7300 12004 7306 12006
rect 8201 12003 8267 12006
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 3141 11932 3207 11933
rect 2814 11930 2820 11932
rect 0 11870 2820 11930
rect 0 11840 800 11870
rect 2814 11868 2820 11870
rect 2884 11868 2890 11932
rect 3141 11928 3188 11932
rect 3252 11930 3258 11932
rect 22200 11930 23000 11960
rect 3141 11872 3146 11928
rect 3141 11868 3188 11872
rect 3252 11870 3298 11930
rect 3252 11868 3258 11870
rect 3141 11867 3207 11868
rect 22142 11840 23000 11930
rect 2313 11794 2379 11797
rect 10133 11794 10199 11797
rect 18045 11794 18111 11797
rect 22142 11794 22202 11840
rect 2313 11792 12450 11794
rect 2313 11736 2318 11792
rect 2374 11736 10138 11792
rect 10194 11736 12450 11792
rect 2313 11734 12450 11736
rect 2313 11731 2379 11734
rect 10133 11731 10199 11734
rect 12390 11658 12450 11734
rect 18045 11792 22202 11794
rect 18045 11736 18050 11792
rect 18106 11736 22202 11792
rect 18045 11734 22202 11736
rect 18045 11731 18111 11734
rect 14273 11658 14339 11661
rect 12390 11656 14339 11658
rect 12390 11600 14278 11656
rect 14334 11600 14339 11656
rect 12390 11598 14339 11600
rect 14273 11595 14339 11598
rect 18597 11658 18663 11661
rect 18597 11656 19626 11658
rect 18597 11600 18602 11656
rect 18658 11600 19626 11656
rect 18597 11598 19626 11600
rect 18597 11595 18663 11598
rect 0 11522 800 11552
rect 3049 11522 3115 11525
rect 0 11520 3115 11522
rect 0 11464 3054 11520
rect 3110 11464 3115 11520
rect 0 11462 3115 11464
rect 19566 11522 19626 11598
rect 22200 11522 23000 11552
rect 19566 11462 23000 11522
rect 0 11432 800 11462
rect 3049 11459 3115 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 0 11114 800 11144
rect 3366 11114 3372 11116
rect 0 11054 3372 11114
rect 0 11024 800 11054
rect 3366 11052 3372 11054
rect 3436 11052 3442 11116
rect 4337 11114 4403 11117
rect 4470 11114 4476 11116
rect 4337 11112 4476 11114
rect 4337 11056 4342 11112
rect 4398 11056 4476 11112
rect 4337 11054 4476 11056
rect 4337 11051 4403 11054
rect 4470 11052 4476 11054
rect 4540 11052 4546 11116
rect 6913 11114 6979 11117
rect 14641 11114 14707 11117
rect 6913 11112 14707 11114
rect 6913 11056 6918 11112
rect 6974 11056 14646 11112
rect 14702 11056 14707 11112
rect 6913 11054 14707 11056
rect 6913 11051 6979 11054
rect 14641 11051 14707 11054
rect 20253 11114 20319 11117
rect 22200 11114 23000 11144
rect 20253 11112 23000 11114
rect 20253 11056 20258 11112
rect 20314 11056 23000 11112
rect 20253 11054 23000 11056
rect 20253 11051 20319 11054
rect 22200 11024 23000 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 7741 10842 7807 10845
rect 7925 10842 7991 10845
rect 7741 10840 7991 10842
rect 7741 10784 7746 10840
rect 7802 10784 7930 10840
rect 7986 10784 7991 10840
rect 7741 10782 7991 10784
rect 7741 10779 7807 10782
rect 7925 10779 7991 10782
rect 0 10706 800 10736
rect 4889 10706 4955 10709
rect 10174 10706 10180 10708
rect 0 10646 3986 10706
rect 0 10616 800 10646
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 3926 10298 3986 10646
rect 4889 10704 10180 10706
rect 4889 10648 4894 10704
rect 4950 10648 10180 10704
rect 4889 10646 10180 10648
rect 4889 10643 4955 10646
rect 10174 10644 10180 10646
rect 10244 10706 10250 10708
rect 22200 10706 23000 10736
rect 10244 10646 23000 10706
rect 10244 10644 10250 10646
rect 22200 10616 23000 10646
rect 4061 10570 4127 10573
rect 10685 10570 10751 10573
rect 4061 10568 10751 10570
rect 4061 10512 4066 10568
rect 4122 10512 10690 10568
rect 10746 10512 10751 10568
rect 4061 10510 10751 10512
rect 4061 10507 4127 10510
rect 10685 10507 10751 10510
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 22200 10298 23000 10328
rect 0 10238 2146 10298
rect 3926 10238 4124 10298
rect 0 10208 800 10238
rect 2086 10162 2146 10238
rect 3877 10162 3943 10165
rect 2086 10160 3943 10162
rect 2086 10104 3882 10160
rect 3938 10104 3943 10160
rect 2086 10102 3943 10104
rect 4064 10162 4124 10238
rect 19566 10238 23000 10298
rect 11094 10162 11100 10164
rect 4064 10102 11100 10162
rect 3877 10099 3943 10102
rect 11094 10100 11100 10102
rect 11164 10100 11170 10164
rect 12157 10162 12223 10165
rect 19566 10162 19626 10238
rect 22200 10208 23000 10238
rect 12157 10160 19626 10162
rect 12157 10104 12162 10160
rect 12218 10104 19626 10160
rect 12157 10102 19626 10104
rect 12157 10099 12223 10102
rect 6085 10026 6151 10029
rect 7925 10026 7991 10029
rect 10593 10026 10659 10029
rect 6085 10024 10659 10026
rect 6085 9968 6090 10024
rect 6146 9968 7930 10024
rect 7986 9968 10598 10024
rect 10654 9968 10659 10024
rect 6085 9966 10659 9968
rect 6085 9963 6151 9966
rect 7925 9963 7991 9966
rect 10593 9963 10659 9966
rect 17953 10026 18019 10029
rect 17953 10024 22202 10026
rect 17953 9968 17958 10024
rect 18014 9968 22202 10024
rect 17953 9966 22202 9968
rect 17953 9963 18019 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 4061 9890 4127 9893
rect 0 9888 4127 9890
rect 0 9832 4066 9888
rect 4122 9832 4127 9888
rect 0 9830 4127 9832
rect 0 9800 800 9830
rect 4061 9827 4127 9830
rect 19425 9890 19491 9893
rect 19558 9890 19564 9892
rect 19425 9888 19564 9890
rect 19425 9832 19430 9888
rect 19486 9832 19564 9888
rect 19425 9830 19564 9832
rect 19425 9827 19491 9830
rect 19558 9828 19564 9830
rect 19628 9828 19634 9892
rect 22142 9830 23000 9920
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 3601 9618 3667 9621
rect 5206 9618 5212 9620
rect 3601 9616 5212 9618
rect 3601 9560 3606 9616
rect 3662 9560 5212 9616
rect 3601 9558 5212 9560
rect 3601 9555 3667 9558
rect 5206 9556 5212 9558
rect 5276 9556 5282 9620
rect 0 9482 800 9512
rect 4153 9482 4219 9485
rect 0 9480 4219 9482
rect 0 9424 4158 9480
rect 4214 9424 4219 9480
rect 0 9422 4219 9424
rect 0 9392 800 9422
rect 4153 9419 4219 9422
rect 4705 9482 4771 9485
rect 9029 9482 9095 9485
rect 4705 9480 9095 9482
rect 4705 9424 4710 9480
rect 4766 9424 9034 9480
rect 9090 9424 9095 9480
rect 4705 9422 9095 9424
rect 4705 9419 4771 9422
rect 9029 9419 9095 9422
rect 18597 9482 18663 9485
rect 22200 9482 23000 9512
rect 18597 9480 23000 9482
rect 18597 9424 18602 9480
rect 18658 9424 23000 9480
rect 18597 9422 23000 9424
rect 18597 9419 18663 9422
rect 22200 9392 23000 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 3325 9210 3391 9213
rect 2730 9208 3391 9210
rect 2730 9152 3330 9208
rect 3386 9152 3391 9208
rect 2730 9150 3391 9152
rect 0 9074 800 9104
rect 2730 9074 2790 9150
rect 3325 9147 3391 9150
rect 0 9014 2790 9074
rect 17953 9074 18019 9077
rect 22200 9074 23000 9104
rect 17953 9072 23000 9074
rect 17953 9016 17958 9072
rect 18014 9016 23000 9072
rect 17953 9014 23000 9016
rect 0 8984 800 9014
rect 17953 9011 18019 9014
rect 22200 8984 23000 9014
rect 8201 8938 8267 8941
rect 12249 8938 12315 8941
rect 8201 8936 12315 8938
rect 8201 8880 8206 8936
rect 8262 8880 12254 8936
rect 12310 8880 12315 8936
rect 8201 8878 12315 8880
rect 8201 8875 8267 8878
rect 12249 8875 12315 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 4061 8666 4127 8669
rect 22200 8666 23000 8696
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 800 8606
rect 4061 8603 4127 8606
rect 22142 8576 23000 8666
rect 18137 8530 18203 8533
rect 22142 8530 22202 8576
rect 18137 8528 22202 8530
rect 18137 8472 18142 8528
rect 18198 8472 22202 8528
rect 18137 8470 22202 8472
rect 18137 8467 18203 8470
rect 4102 8332 4108 8396
rect 4172 8394 4178 8396
rect 4245 8394 4311 8397
rect 4172 8392 4311 8394
rect 4172 8336 4250 8392
rect 4306 8336 4311 8392
rect 4172 8334 4311 8336
rect 4172 8332 4178 8334
rect 4245 8331 4311 8334
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 10317 8258 10383 8261
rect 13077 8258 13143 8261
rect 22200 8258 23000 8288
rect 10317 8256 13143 8258
rect 10317 8200 10322 8256
rect 10378 8200 13082 8256
rect 13138 8200 13143 8256
rect 10317 8198 13143 8200
rect 10317 8195 10383 8198
rect 13077 8195 13143 8198
rect 19566 8198 23000 8258
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 6678 8060 6684 8124
rect 6748 8122 6754 8124
rect 7649 8122 7715 8125
rect 6748 8120 7715 8122
rect 6748 8064 7654 8120
rect 7710 8064 7715 8120
rect 6748 8062 7715 8064
rect 6748 8060 6754 8062
rect 7649 8059 7715 8062
rect 9857 7986 9923 7989
rect 19566 7986 19626 8198
rect 22200 8168 23000 8198
rect 9857 7984 19626 7986
rect 9857 7928 9862 7984
rect 9918 7928 19626 7984
rect 9857 7926 19626 7928
rect 9857 7923 9923 7926
rect 0 7850 800 7880
rect 1577 7850 1643 7853
rect 0 7848 1643 7850
rect 0 7792 1582 7848
rect 1638 7792 1643 7848
rect 0 7790 1643 7792
rect 0 7760 800 7790
rect 1577 7787 1643 7790
rect 4889 7850 4955 7853
rect 10317 7850 10383 7853
rect 4889 7848 10383 7850
rect 4889 7792 4894 7848
rect 4950 7792 10322 7848
rect 10378 7792 10383 7848
rect 4889 7790 10383 7792
rect 4889 7787 4955 7790
rect 10317 7787 10383 7790
rect 17769 7850 17835 7853
rect 22200 7850 23000 7880
rect 17769 7848 23000 7850
rect 17769 7792 17774 7848
rect 17830 7792 23000 7848
rect 17769 7790 23000 7792
rect 17769 7787 17835 7790
rect 22200 7760 23000 7790
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 3969 7578 4035 7581
rect 2730 7576 4035 7578
rect 2730 7520 3974 7576
rect 4030 7520 4035 7576
rect 2730 7518 4035 7520
rect 0 7442 800 7472
rect 2730 7442 2790 7518
rect 3969 7515 4035 7518
rect 5441 7442 5507 7445
rect 17493 7442 17559 7445
rect 0 7382 2790 7442
rect 3374 7440 17559 7442
rect 3374 7384 5446 7440
rect 5502 7384 17498 7440
rect 17554 7384 17559 7440
rect 3374 7382 17559 7384
rect 0 7352 800 7382
rect 0 7034 800 7064
rect 3374 7034 3434 7382
rect 5441 7379 5507 7382
rect 17493 7379 17559 7382
rect 18045 7442 18111 7445
rect 22200 7442 23000 7472
rect 18045 7440 23000 7442
rect 18045 7384 18050 7440
rect 18106 7384 23000 7440
rect 18045 7382 23000 7384
rect 18045 7379 18111 7382
rect 22200 7352 23000 7382
rect 6821 7306 6887 7309
rect 9305 7306 9371 7309
rect 10961 7306 11027 7309
rect 6821 7304 11027 7306
rect 6821 7248 6826 7304
rect 6882 7248 9310 7304
rect 9366 7248 10966 7304
rect 11022 7248 11027 7304
rect 6821 7246 11027 7248
rect 6821 7243 6887 7246
rect 9305 7243 9371 7246
rect 10961 7243 11027 7246
rect 18229 7306 18295 7309
rect 18229 7304 20730 7306
rect 18229 7248 18234 7304
rect 18290 7248 20730 7304
rect 18229 7246 20730 7248
rect 18229 7243 18295 7246
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 20529 7034 20595 7037
rect 0 6974 3434 7034
rect 20486 7032 20595 7034
rect 20486 6976 20534 7032
rect 20590 6976 20595 7032
rect 0 6944 800 6974
rect 20486 6971 20595 6976
rect 20670 7034 20730 7246
rect 22200 7034 23000 7064
rect 20670 6974 23000 7034
rect 4521 6900 4587 6901
rect 4470 6898 4476 6900
rect 4430 6838 4476 6898
rect 4540 6898 4587 6900
rect 9581 6898 9647 6901
rect 4540 6896 9647 6898
rect 4582 6840 9586 6896
rect 9642 6840 9647 6896
rect 4470 6836 4476 6838
rect 4540 6838 9647 6840
rect 4540 6836 4587 6838
rect 4521 6835 4587 6836
rect 9581 6835 9647 6838
rect 7046 6700 7052 6764
rect 7116 6762 7122 6764
rect 18781 6762 18847 6765
rect 20486 6762 20546 6971
rect 22200 6944 23000 6974
rect 7116 6760 20546 6762
rect 7116 6704 18786 6760
rect 18842 6704 20546 6760
rect 7116 6702 20546 6704
rect 20670 6702 22202 6762
rect 7116 6700 7122 6702
rect 18781 6699 18847 6702
rect 0 6626 800 6656
rect 3141 6628 3207 6629
rect 3141 6626 3188 6628
rect 0 6566 2790 6626
rect 3096 6624 3188 6626
rect 3096 6568 3146 6624
rect 3096 6566 3188 6568
rect 0 6536 800 6566
rect 2730 6490 2790 6566
rect 3141 6564 3188 6566
rect 3252 6564 3258 6628
rect 17677 6626 17743 6629
rect 20670 6626 20730 6702
rect 17677 6624 20730 6626
rect 17677 6568 17682 6624
rect 17738 6568 20730 6624
rect 17677 6566 20730 6568
rect 22142 6656 22202 6702
rect 22142 6566 23000 6656
rect 3141 6563 3207 6564
rect 17677 6563 17743 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 4061 6490 4127 6493
rect 2730 6488 4127 6490
rect 2730 6432 4066 6488
rect 4122 6432 4127 6488
rect 2730 6430 4127 6432
rect 4061 6427 4127 6430
rect 3969 6354 4035 6357
rect 8845 6354 8911 6357
rect 3969 6352 8911 6354
rect 3969 6296 3974 6352
rect 4030 6296 8850 6352
rect 8906 6296 8911 6352
rect 3969 6294 8911 6296
rect 3969 6291 4035 6294
rect 8845 6291 8911 6294
rect 9581 6354 9647 6357
rect 15929 6354 15995 6357
rect 9581 6352 15995 6354
rect 9581 6296 9586 6352
rect 9642 6296 15934 6352
rect 15990 6296 15995 6352
rect 9581 6294 15995 6296
rect 9581 6291 9647 6294
rect 15929 6291 15995 6294
rect 0 6218 800 6248
rect 3785 6218 3851 6221
rect 0 6216 3851 6218
rect 0 6160 3790 6216
rect 3846 6160 3851 6216
rect 0 6158 3851 6160
rect 0 6128 800 6158
rect 3785 6155 3851 6158
rect 3969 6218 4035 6221
rect 8753 6218 8819 6221
rect 3969 6216 8819 6218
rect 3969 6160 3974 6216
rect 4030 6160 8758 6216
rect 8814 6160 8819 6216
rect 3969 6158 8819 6160
rect 3969 6155 4035 6158
rect 8753 6155 8819 6158
rect 8937 6218 9003 6221
rect 17033 6218 17099 6221
rect 8937 6216 17099 6218
rect 8937 6160 8942 6216
rect 8998 6160 17038 6216
rect 17094 6160 17099 6216
rect 8937 6158 17099 6160
rect 8937 6155 9003 6158
rect 17033 6155 17099 6158
rect 18505 6218 18571 6221
rect 22200 6218 23000 6248
rect 18505 6216 23000 6218
rect 18505 6160 18510 6216
rect 18566 6160 23000 6216
rect 18505 6158 23000 6160
rect 18505 6155 18571 6158
rect 22200 6128 23000 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 0 5810 800 5840
rect 2814 5810 2820 5812
rect 0 5750 2820 5810
rect 0 5720 800 5750
rect 2814 5748 2820 5750
rect 2884 5748 2890 5812
rect 17902 5748 17908 5812
rect 17972 5810 17978 5812
rect 22200 5810 23000 5840
rect 17972 5750 23000 5810
rect 17972 5748 17978 5750
rect 22200 5720 23000 5750
rect 5717 5674 5783 5677
rect 6453 5674 6519 5677
rect 9305 5674 9371 5677
rect 5717 5672 9371 5674
rect 5717 5616 5722 5672
rect 5778 5616 6458 5672
rect 6514 5616 9310 5672
rect 9366 5616 9371 5672
rect 5717 5614 9371 5616
rect 5717 5611 5783 5614
rect 6453 5611 6519 5614
rect 9305 5611 9371 5614
rect 9673 5674 9739 5677
rect 17309 5674 17375 5677
rect 9673 5672 17375 5674
rect 9673 5616 9678 5672
rect 9734 5616 17314 5672
rect 17370 5616 17375 5672
rect 9673 5614 17375 5616
rect 9673 5611 9739 5614
rect 17309 5611 17375 5614
rect 2589 5538 2655 5541
rect 4102 5538 4108 5540
rect 2589 5536 4108 5538
rect 2589 5480 2594 5536
rect 2650 5480 4108 5536
rect 2589 5478 4108 5480
rect 2589 5475 2655 5478
rect 4102 5476 4108 5478
rect 4172 5476 4178 5540
rect 8017 5538 8083 5541
rect 8150 5538 8156 5540
rect 8017 5536 8156 5538
rect 8017 5480 8022 5536
rect 8078 5480 8156 5536
rect 8017 5478 8156 5480
rect 8017 5475 8083 5478
rect 8150 5476 8156 5478
rect 8220 5476 8226 5540
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 2129 5402 2195 5405
rect 3049 5402 3115 5405
rect 0 5400 3115 5402
rect 0 5344 2134 5400
rect 2190 5344 3054 5400
rect 3110 5344 3115 5400
rect 0 5342 3115 5344
rect 0 5312 800 5342
rect 2129 5339 2195 5342
rect 3049 5339 3115 5342
rect 6637 5402 6703 5405
rect 11053 5402 11119 5405
rect 22200 5402 23000 5432
rect 6637 5400 11119 5402
rect 6637 5344 6642 5400
rect 6698 5344 11058 5400
rect 11114 5344 11119 5400
rect 6637 5342 11119 5344
rect 6637 5339 6703 5342
rect 11053 5339 11119 5342
rect 22142 5312 23000 5402
rect 16573 5266 16639 5269
rect 18505 5266 18571 5269
rect 16573 5264 18571 5266
rect 16573 5208 16578 5264
rect 16634 5208 18510 5264
rect 18566 5208 18571 5264
rect 16573 5206 18571 5208
rect 16573 5203 16639 5206
rect 18505 5203 18571 5206
rect 21265 5266 21331 5269
rect 22142 5266 22202 5312
rect 21265 5264 22202 5266
rect 21265 5208 21270 5264
rect 21326 5208 22202 5264
rect 21265 5206 22202 5208
rect 21265 5203 21331 5206
rect 20529 5132 20595 5133
rect 20478 5068 20484 5132
rect 20548 5130 20595 5132
rect 20548 5128 20640 5130
rect 20590 5072 20640 5128
rect 20548 5070 20640 5072
rect 20548 5068 20595 5070
rect 20529 5067 20595 5068
rect 0 4994 800 5024
rect 1945 4994 2011 4997
rect 0 4992 2011 4994
rect 0 4936 1950 4992
rect 2006 4936 2011 4992
rect 0 4934 2011 4936
rect 0 4904 800 4934
rect 1945 4931 2011 4934
rect 20253 4994 20319 4997
rect 22200 4994 23000 5024
rect 20253 4992 23000 4994
rect 20253 4936 20258 4992
rect 20314 4936 23000 4992
rect 20253 4934 23000 4936
rect 20253 4931 20319 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 4061 4722 4127 4725
rect 10777 4722 10843 4725
rect 4061 4720 10843 4722
rect 4061 4664 4066 4720
rect 4122 4664 10782 4720
rect 10838 4664 10843 4720
rect 4061 4662 10843 4664
rect 4061 4659 4127 4662
rect 10777 4659 10843 4662
rect 0 4586 800 4616
rect 2773 4586 2839 4589
rect 0 4584 2839 4586
rect 0 4528 2778 4584
rect 2834 4528 2839 4584
rect 0 4526 2839 4528
rect 0 4496 800 4526
rect 2773 4523 2839 4526
rect 4429 4586 4495 4589
rect 7230 4586 7236 4588
rect 4429 4584 7236 4586
rect 4429 4528 4434 4584
rect 4490 4528 7236 4584
rect 4429 4526 7236 4528
rect 4429 4523 4495 4526
rect 7230 4524 7236 4526
rect 7300 4586 7306 4588
rect 17902 4586 17908 4588
rect 7300 4526 17908 4586
rect 7300 4524 7306 4526
rect 17902 4524 17908 4526
rect 17972 4524 17978 4588
rect 21173 4586 21239 4589
rect 22200 4586 23000 4616
rect 21173 4584 23000 4586
rect 21173 4528 21178 4584
rect 21234 4528 23000 4584
rect 21173 4526 23000 4528
rect 21173 4523 21239 4526
rect 22200 4496 23000 4526
rect 18597 4450 18663 4453
rect 20989 4450 21055 4453
rect 18597 4448 21055 4450
rect 18597 4392 18602 4448
rect 18658 4392 20994 4448
rect 21050 4392 21055 4448
rect 18597 4390 21055 4392
rect 18597 4387 18663 4390
rect 20989 4387 21055 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 15377 4314 15443 4317
rect 21265 4314 21331 4317
rect 11838 4312 15443 4314
rect 11838 4256 15382 4312
rect 15438 4256 15443 4312
rect 11838 4254 15443 4256
rect 0 4178 800 4208
rect 2865 4178 2931 4181
rect 0 4176 2931 4178
rect 0 4120 2870 4176
rect 2926 4120 2931 4176
rect 0 4118 2931 4120
rect 0 4088 800 4118
rect 2865 4115 2931 4118
rect 5165 4178 5231 4181
rect 8937 4178 9003 4181
rect 5165 4176 9003 4178
rect 5165 4120 5170 4176
rect 5226 4120 8942 4176
rect 8998 4120 9003 4176
rect 5165 4118 9003 4120
rect 5165 4115 5231 4118
rect 8937 4115 9003 4118
rect 9397 4178 9463 4181
rect 11838 4178 11898 4254
rect 15377 4251 15443 4254
rect 17542 4312 21331 4314
rect 17542 4256 21270 4312
rect 21326 4256 21331 4312
rect 17542 4254 21331 4256
rect 9397 4176 11898 4178
rect 9397 4120 9402 4176
rect 9458 4120 11898 4176
rect 9397 4118 11898 4120
rect 13077 4178 13143 4181
rect 17542 4178 17602 4254
rect 21265 4251 21331 4254
rect 13077 4176 17602 4178
rect 13077 4120 13082 4176
rect 13138 4120 17602 4176
rect 13077 4118 17602 4120
rect 17769 4178 17835 4181
rect 19977 4178 20043 4181
rect 17769 4176 20043 4178
rect 17769 4120 17774 4176
rect 17830 4120 19982 4176
rect 20038 4120 20043 4176
rect 17769 4118 20043 4120
rect 9397 4115 9463 4118
rect 13077 4115 13143 4118
rect 17769 4115 17835 4118
rect 19977 4115 20043 4118
rect 20989 4178 21055 4181
rect 22200 4178 23000 4208
rect 20989 4176 23000 4178
rect 20989 4120 20994 4176
rect 21050 4120 23000 4176
rect 20989 4118 23000 4120
rect 20989 4115 21055 4118
rect 22200 4088 23000 4118
rect 2129 4042 2195 4045
rect 2814 4042 2820 4044
rect 2129 4040 2820 4042
rect 2129 3984 2134 4040
rect 2190 3984 2820 4040
rect 2129 3982 2820 3984
rect 2129 3979 2195 3982
rect 2814 3980 2820 3982
rect 2884 4042 2890 4044
rect 7925 4042 7991 4045
rect 2884 4040 7991 4042
rect 2884 3984 7930 4040
rect 7986 3984 7991 4040
rect 2884 3982 7991 3984
rect 2884 3980 2890 3982
rect 7925 3979 7991 3982
rect 9305 4042 9371 4045
rect 9438 4042 9444 4044
rect 9305 4040 9444 4042
rect 9305 3984 9310 4040
rect 9366 3984 9444 4040
rect 9305 3982 9444 3984
rect 9305 3979 9371 3982
rect 9438 3980 9444 3982
rect 9508 3980 9514 4044
rect 9581 4042 9647 4045
rect 18413 4042 18479 4045
rect 19333 4042 19399 4045
rect 9581 4040 19399 4042
rect 9581 3984 9586 4040
rect 9642 3984 18418 4040
rect 18474 3984 19338 4040
rect 19394 3984 19399 4040
rect 9581 3982 19399 3984
rect 9581 3979 9647 3982
rect 18413 3979 18479 3982
rect 19333 3979 19399 3982
rect 9806 3844 9812 3908
rect 9876 3906 9882 3908
rect 10685 3906 10751 3909
rect 9876 3904 10751 3906
rect 9876 3848 10690 3904
rect 10746 3848 10751 3904
rect 9876 3846 10751 3848
rect 9876 3844 9882 3846
rect 10685 3843 10751 3846
rect 11145 3906 11211 3909
rect 11329 3906 11395 3909
rect 11145 3904 11395 3906
rect 11145 3848 11150 3904
rect 11206 3848 11334 3904
rect 11390 3848 11395 3904
rect 11145 3846 11395 3848
rect 11145 3843 11211 3846
rect 11329 3843 11395 3846
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 1393 3770 1459 3773
rect 13813 3770 13879 3773
rect 0 3768 1459 3770
rect 0 3712 1398 3768
rect 1454 3712 1459 3768
rect 0 3710 1459 3712
rect 0 3680 800 3710
rect 1393 3707 1459 3710
rect 9262 3768 13879 3770
rect 9262 3712 13818 3768
rect 13874 3712 13879 3768
rect 9262 3710 13879 3712
rect 5533 3634 5599 3637
rect 9262 3634 9322 3710
rect 13813 3707 13879 3710
rect 21357 3770 21423 3773
rect 22200 3770 23000 3800
rect 21357 3768 23000 3770
rect 21357 3712 21362 3768
rect 21418 3712 23000 3768
rect 21357 3710 23000 3712
rect 21357 3707 21423 3710
rect 22200 3680 23000 3710
rect 13261 3634 13327 3637
rect 5533 3632 9322 3634
rect 5533 3576 5538 3632
rect 5594 3576 9322 3632
rect 5533 3574 9322 3576
rect 9630 3632 13327 3634
rect 9630 3576 13266 3632
rect 13322 3576 13327 3632
rect 9630 3574 13327 3576
rect 5533 3571 5599 3574
rect 5758 3436 5764 3500
rect 5828 3498 5834 3500
rect 8937 3498 9003 3501
rect 5828 3496 9003 3498
rect 5828 3440 8942 3496
rect 8998 3440 9003 3496
rect 5828 3438 9003 3440
rect 5828 3436 5834 3438
rect 8937 3435 9003 3438
rect 0 3362 800 3392
rect 1761 3362 1827 3365
rect 7005 3364 7071 3365
rect 9213 3364 9279 3365
rect 7005 3362 7052 3364
rect 0 3360 1827 3362
rect 0 3304 1766 3360
rect 1822 3304 1827 3360
rect 0 3302 1827 3304
rect 6960 3360 7052 3362
rect 6960 3304 7010 3360
rect 6960 3302 7052 3304
rect 0 3272 800 3302
rect 1761 3299 1827 3302
rect 7005 3300 7052 3302
rect 7116 3300 7122 3364
rect 9213 3360 9260 3364
rect 9324 3362 9330 3364
rect 9213 3304 9218 3360
rect 9213 3300 9260 3304
rect 9324 3302 9370 3362
rect 9324 3300 9330 3302
rect 7005 3299 7071 3300
rect 9213 3299 9279 3300
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 6729 3226 6795 3229
rect 9630 3226 9690 3574
rect 13261 3571 13327 3574
rect 16665 3634 16731 3637
rect 18321 3634 18387 3637
rect 16665 3632 18387 3634
rect 16665 3576 16670 3632
rect 16726 3576 18326 3632
rect 18382 3576 18387 3632
rect 16665 3574 18387 3576
rect 16665 3571 16731 3574
rect 18321 3571 18387 3574
rect 18965 3498 19031 3501
rect 21449 3498 21515 3501
rect 18965 3496 22202 3498
rect 18965 3440 18970 3496
rect 19026 3440 21454 3496
rect 21510 3440 22202 3496
rect 18965 3438 22202 3440
rect 18965 3435 19031 3438
rect 21449 3435 21515 3438
rect 22142 3392 22202 3438
rect 22142 3302 23000 3392
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 6729 3224 9690 3226
rect 6729 3168 6734 3224
rect 6790 3168 9690 3224
rect 6729 3166 9690 3168
rect 6729 3163 6795 3166
rect 5809 3090 5875 3093
rect 14457 3090 14523 3093
rect 5809 3088 14523 3090
rect 5809 3032 5814 3088
rect 5870 3032 14462 3088
rect 14518 3032 14523 3088
rect 5809 3030 14523 3032
rect 5809 3027 5875 3030
rect 14457 3027 14523 3030
rect 0 2954 800 2984
rect 3325 2954 3391 2957
rect 0 2952 3391 2954
rect 0 2896 3330 2952
rect 3386 2896 3391 2952
rect 0 2894 3391 2896
rect 0 2864 800 2894
rect 3325 2891 3391 2894
rect 7741 2954 7807 2957
rect 13813 2954 13879 2957
rect 7741 2952 13879 2954
rect 7741 2896 7746 2952
rect 7802 2896 13818 2952
rect 13874 2896 13879 2952
rect 7741 2894 13879 2896
rect 7741 2891 7807 2894
rect 13813 2891 13879 2894
rect 18505 2954 18571 2957
rect 18873 2954 18939 2957
rect 18505 2952 18939 2954
rect 18505 2896 18510 2952
rect 18566 2896 18878 2952
rect 18934 2896 18939 2952
rect 18505 2894 18939 2896
rect 18505 2891 18571 2894
rect 18873 2891 18939 2894
rect 20805 2954 20871 2957
rect 22200 2954 23000 2984
rect 20805 2952 23000 2954
rect 20805 2896 20810 2952
rect 20866 2896 23000 2952
rect 20805 2894 23000 2896
rect 20805 2891 20871 2894
rect 22200 2864 23000 2894
rect 9765 2818 9831 2821
rect 10225 2818 10291 2821
rect 9765 2816 10291 2818
rect 9765 2760 9770 2816
rect 9826 2760 10230 2816
rect 10286 2760 10291 2816
rect 9765 2758 10291 2760
rect 9765 2755 9831 2758
rect 10225 2755 10291 2758
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 0 2546 800 2576
rect 3233 2546 3299 2549
rect 0 2544 3299 2546
rect 0 2488 3238 2544
rect 3294 2488 3299 2544
rect 0 2486 3299 2488
rect 0 2456 800 2486
rect 3233 2483 3299 2486
rect 6913 2546 6979 2549
rect 9622 2546 9628 2548
rect 6913 2544 9628 2546
rect 6913 2488 6918 2544
rect 6974 2488 9628 2544
rect 6913 2486 9628 2488
rect 6913 2483 6979 2486
rect 9622 2484 9628 2486
rect 9692 2484 9698 2548
rect 18965 2546 19031 2549
rect 20989 2546 21055 2549
rect 22200 2546 23000 2576
rect 18965 2544 23000 2546
rect 18965 2488 18970 2544
rect 19026 2488 20994 2544
rect 21050 2488 23000 2544
rect 18965 2486 23000 2488
rect 18965 2483 19031 2486
rect 20989 2483 21055 2486
rect 22200 2456 23000 2486
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 1853 2138 1919 2141
rect 22200 2138 23000 2168
rect 0 2136 1919 2138
rect 0 2080 1858 2136
rect 1914 2080 1919 2136
rect 0 2078 1919 2080
rect 0 2048 800 2078
rect 1853 2075 1919 2078
rect 22142 2048 23000 2138
rect 21081 2002 21147 2005
rect 22142 2002 22202 2048
rect 21081 2000 22202 2002
rect 21081 1944 21086 2000
rect 21142 1944 22202 2000
rect 21081 1942 22202 1944
rect 21081 1939 21147 1942
rect 0 1730 800 1760
rect 3417 1730 3483 1733
rect 0 1728 3483 1730
rect 0 1672 3422 1728
rect 3478 1672 3483 1728
rect 0 1670 3483 1672
rect 0 1640 800 1670
rect 3417 1667 3483 1670
rect 18689 1730 18755 1733
rect 22200 1730 23000 1760
rect 18689 1728 23000 1730
rect 18689 1672 18694 1728
rect 18750 1672 23000 1728
rect 18689 1670 23000 1672
rect 18689 1667 18755 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 11100 19680 11164 19684
rect 11100 19624 11114 19680
rect 11114 19624 11164 19680
rect 11100 19620 11164 19624
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3372 19348 3436 19412
rect 9260 19348 9324 19412
rect 16988 19348 17052 19412
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 19564 18124 19628 18188
rect 5212 17988 5276 18052
rect 10180 18048 10244 18052
rect 10180 17992 10194 18048
rect 10194 17992 10244 18048
rect 10180 17988 10244 17992
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 10548 17036 10612 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 4292 16628 4356 16692
rect 6684 16628 6748 16692
rect 8156 16628 8220 16692
rect 20484 16628 20548 16692
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 7052 15948 7116 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 9444 15404 9508 15468
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 16988 14996 17052 15060
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 2820 13364 2884 13428
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 9628 13364 9692 13428
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 8340 12820 8404 12884
rect 10548 12684 10612 12748
rect 5764 12548 5828 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 4292 12276 4356 12340
rect 4476 12276 4540 12340
rect 8340 12276 8404 12340
rect 9812 12276 9876 12340
rect 7236 12004 7300 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 2820 11868 2884 11932
rect 3188 11928 3252 11932
rect 3188 11872 3202 11928
rect 3202 11872 3252 11928
rect 3188 11868 3252 11872
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 3372 11052 3436 11116
rect 4476 11052 4540 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 10180 10644 10244 10708
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 11100 10100 11164 10164
rect 19564 9828 19628 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 5212 9556 5276 9620
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 4108 8332 4172 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6684 8060 6748 8124
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 4476 6896 4540 6900
rect 4476 6840 4526 6896
rect 4526 6840 4540 6896
rect 4476 6836 4540 6840
rect 7052 6700 7116 6764
rect 3188 6624 3252 6628
rect 3188 6568 3202 6624
rect 3202 6568 3252 6624
rect 3188 6564 3252 6568
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 2820 5748 2884 5812
rect 17908 5748 17972 5812
rect 4108 5476 4172 5540
rect 8156 5476 8220 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 20484 5128 20548 5132
rect 20484 5072 20534 5128
rect 20534 5072 20548 5128
rect 20484 5068 20548 5072
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 7236 4524 7300 4588
rect 17908 4524 17972 4588
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 2820 3980 2884 4044
rect 9444 3980 9508 4044
rect 9812 3844 9876 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 5764 3436 5828 3500
rect 7052 3360 7116 3364
rect 7052 3304 7066 3360
rect 7066 3304 7116 3360
rect 7052 3300 7116 3304
rect 9260 3360 9324 3364
rect 9260 3304 9274 3360
rect 9274 3304 9324 3360
rect 9260 3300 9324 3304
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 9628 2484 9692 2548
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3371 19412 3437 19413
rect 3371 19348 3372 19412
rect 3436 19348 3437 19412
rect 3371 19347 3437 19348
rect 2819 13428 2885 13429
rect 2819 13364 2820 13428
rect 2884 13364 2885 13428
rect 2819 13363 2885 13364
rect 2822 11933 2882 13363
rect 2819 11932 2885 11933
rect 2819 11868 2820 11932
rect 2884 11868 2885 11932
rect 2819 11867 2885 11868
rect 3187 11932 3253 11933
rect 3187 11868 3188 11932
rect 3252 11868 3253 11932
rect 3187 11867 3253 11868
rect 3190 6629 3250 11867
rect 3374 11117 3434 19347
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5211 18052 5277 18053
rect 5211 17988 5212 18052
rect 5276 17988 5277 18052
rect 5211 17987 5277 17988
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 4291 16692 4357 16693
rect 4291 16628 4292 16692
rect 4356 16628 4357 16692
rect 4291 16627 4357 16628
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 4294 12341 4354 16627
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 4475 12340 4541 12341
rect 4475 12276 4476 12340
rect 4540 12276 4541 12340
rect 4475 12275 4541 12276
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 3543 10368 3863 11392
rect 4478 11117 4538 12275
rect 4475 11116 4541 11117
rect 4475 11052 4476 11116
rect 4540 11052 4541 11116
rect 4475 11051 4541 11052
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 4107 8396 4173 8397
rect 4107 8332 4108 8396
rect 4172 8332 4173 8396
rect 4107 8331 4173 8332
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3187 6628 3253 6629
rect 3187 6564 3188 6628
rect 3252 6564 3253 6628
rect 3187 6563 3253 6564
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 2819 5812 2885 5813
rect 2819 5748 2820 5812
rect 2884 5748 2885 5812
rect 2819 5747 2885 5748
rect 2822 4045 2882 5747
rect 3543 4928 3863 5952
rect 4110 5541 4170 8331
rect 4478 6901 4538 11051
rect 5214 9621 5274 17987
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11099 19684 11165 19685
rect 11099 19620 11100 19684
rect 11164 19620 11165 19684
rect 11099 19619 11165 19620
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 6683 16692 6749 16693
rect 6683 16628 6684 16692
rect 6748 16628 6749 16692
rect 6683 16627 6749 16628
rect 8155 16692 8221 16693
rect 8155 16628 8156 16692
rect 8220 16628 8221 16692
rect 8155 16627 8221 16628
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5763 12612 5829 12613
rect 5763 12548 5764 12612
rect 5828 12548 5829 12612
rect 5763 12547 5829 12548
rect 5211 9620 5277 9621
rect 5211 9556 5212 9620
rect 5276 9556 5277 9620
rect 5211 9555 5277 9556
rect 4475 6900 4541 6901
rect 4475 6836 4476 6900
rect 4540 6836 4541 6900
rect 4475 6835 4541 6836
rect 4107 5540 4173 5541
rect 4107 5476 4108 5540
rect 4172 5476 4173 5540
rect 4107 5475 4173 5476
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 2819 4044 2885 4045
rect 2819 3980 2820 4044
rect 2884 3980 2885 4044
rect 2819 3979 2885 3980
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 5766 3501 5826 12547
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6686 8125 6746 16627
rect 7051 16012 7117 16013
rect 7051 15948 7052 16012
rect 7116 15948 7117 16012
rect 7051 15947 7117 15948
rect 6683 8124 6749 8125
rect 6683 8060 6684 8124
rect 6748 8060 6749 8124
rect 6683 8059 6749 8060
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 7054 6765 7114 15947
rect 7235 12068 7301 12069
rect 7235 12004 7236 12068
rect 7300 12004 7301 12068
rect 7235 12003 7301 12004
rect 7051 6764 7117 6765
rect 7051 6700 7052 6764
rect 7116 6700 7117 6764
rect 7051 6699 7117 6700
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5763 3500 5829 3501
rect 5763 3436 5764 3500
rect 5828 3436 5829 3500
rect 5763 3435 5829 3436
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 7054 3365 7114 6699
rect 7238 4589 7298 12003
rect 8158 5541 8218 16627
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8339 12884 8405 12885
rect 8339 12820 8340 12884
rect 8404 12820 8405 12884
rect 8339 12819 8405 12820
rect 8342 12341 8402 12819
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8339 12340 8405 12341
rect 8339 12276 8340 12340
rect 8404 12276 8405 12340
rect 8339 12275 8405 12276
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8155 5540 8221 5541
rect 8155 5476 8156 5540
rect 8220 5476 8221 5540
rect 8155 5475 8221 5476
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 7235 4588 7301 4589
rect 7235 4524 7236 4588
rect 7300 4524 7301 4588
rect 7235 4523 7301 4524
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7051 3364 7117 3365
rect 7051 3300 7052 3364
rect 7116 3300 7117 3364
rect 7051 3299 7117 3300
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2752 9061 3776
rect 9262 3365 9322 19347
rect 10179 18052 10245 18053
rect 10179 17988 10180 18052
rect 10244 17988 10245 18052
rect 10179 17987 10245 17988
rect 9443 15468 9509 15469
rect 9443 15404 9444 15468
rect 9508 15404 9509 15468
rect 9443 15403 9509 15404
rect 9446 4045 9506 15403
rect 9627 13428 9693 13429
rect 9627 13364 9628 13428
rect 9692 13364 9693 13428
rect 9627 13363 9693 13364
rect 9443 4044 9509 4045
rect 9443 3980 9444 4044
rect 9508 3980 9509 4044
rect 9443 3979 9509 3980
rect 9259 3364 9325 3365
rect 9259 3300 9260 3364
rect 9324 3300 9325 3364
rect 9259 3299 9325 3300
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 9630 2549 9690 13363
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9814 3909 9874 12275
rect 10182 10709 10242 17987
rect 10547 17100 10613 17101
rect 10547 17036 10548 17100
rect 10612 17036 10613 17100
rect 10547 17035 10613 17036
rect 10550 12749 10610 17035
rect 10547 12748 10613 12749
rect 10547 12684 10548 12748
rect 10612 12684 10613 12748
rect 10547 12683 10613 12684
rect 10179 10708 10245 10709
rect 10179 10644 10180 10708
rect 10244 10644 10245 10708
rect 10179 10643 10245 10644
rect 11102 10165 11162 19619
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11099 10164 11165 10165
rect 11099 10100 11100 10164
rect 11164 10100 11165 10164
rect 11099 10099 11165 10100
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 9811 3908 9877 3909
rect 9811 3844 9812 3908
rect 9876 3844 9877 3908
rect 9811 3843 9877 3844
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9627 2548 9693 2549
rect 9627 2484 9628 2548
rect 9692 2484 9693 2548
rect 9627 2483 9693 2484
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 16987 19412 17053 19413
rect 16987 19348 16988 19412
rect 17052 19348 17053 19412
rect 16987 19347 17053 19348
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16990 15061 17050 19347
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 19563 18188 19629 18189
rect 19563 18124 19564 18188
rect 19628 18124 19629 18188
rect 19563 18123 19629 18124
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 16987 15060 17053 15061
rect 16987 14996 16988 15060
rect 17052 14996 17053 15060
rect 16987 14995 17053 14996
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19566 9893 19626 18123
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 20483 16692 20549 16693
rect 20483 16628 20484 16692
rect 20548 16628 20549 16692
rect 20483 16627 20549 16628
rect 19563 9892 19629 9893
rect 19563 9828 19564 9892
rect 19628 9828 19629 9892
rect 19563 9827 19629 9828
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 17907 5812 17973 5813
rect 17907 5748 17908 5812
rect 17972 5748 17973 5812
rect 17907 5747 17973 5748
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 17910 4589 17970 5747
rect 19137 4928 19457 5952
rect 20486 5133 20546 16627
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 20483 5132 20549 5133
rect 20483 5068 20484 5132
rect 20548 5068 20549 5132
rect 20483 5067 20549 5068
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 17907 4588 17973 4589
rect 17907 4524 17908 4588
rect 17972 4524 17973 4588
rect 17907 4523 17973 4524
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1649977179
transform -1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform -1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform -1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform -1 0 1656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 4416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 2576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform -1 0 1656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 2944 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform -1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform -1 0 20424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform -1 0 17112 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 9936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform 1 0 19872 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform -1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform -1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform -1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11592 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17940 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 1472 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 4232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 8096 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 7360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18584 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 6992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6808 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1649977179
transform -1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1649977179
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1649977179
transform 1 0 1472 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 1472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 3404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 9016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1649977179
transform -1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 18676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 12972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1649977179
transform -1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1649977179
transform -1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform -1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1649977179
transform -1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 6716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 7728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 18584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1649977179
transform 1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50
timestamp 1649977179
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_210
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1649977179
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1649977179
transform 1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1649977179
transform 1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1649977179
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1649977179
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_43
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_98
timestamp 1649977179
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1649977179
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1649977179
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_9
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_47
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_63
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_115
timestamp 1649977179
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1649977179
transform 1 0 12144 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_128
timestamp 1649977179
transform 1 0 12880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_139
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_187
timestamp 1649977179
transform 1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_191
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_5
timestamp 1649977179
transform 1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1649977179
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_46
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1649977179
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_10
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1649977179
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_64
timestamp 1649977179
transform 1 0 6992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1649977179
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_122
timestamp 1649977179
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_182
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_186
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_190
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_60
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_74
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_108
timestamp 1649977179
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1649977179
transform 1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_183
timestamp 1649977179
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_187
timestamp 1649977179
transform 1 0 18308 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_25
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_94
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_139
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1649977179
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1649977179
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_5
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_108
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_116
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_143
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_64
timestamp 1649977179
transform 1 0 6992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_68
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_72
timestamp 1649977179
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1649977179
transform 1 0 15824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_35
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_39
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_42
timestamp 1649977179
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_46
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_190
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_30
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_61
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_65
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_71
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_94
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_100
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1649977179
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_171
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1649977179
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_5
timestamp 1649977179
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_23
timestamp 1649977179
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_69
timestamp 1649977179
transform 1 0 7452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_179
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_5
timestamp 1649977179
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_13
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1649977179
transform 1 0 2668 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_61
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_185
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_34
timestamp 1649977179
transform 1 0 4232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1649977179
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_57
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_76
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_124
timestamp 1649977179
transform 1 0 12512 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_158
timestamp 1649977179
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_166
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1649977179
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_208
timestamp 1649977179
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_26
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_30
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1649977179
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_67
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1649977179
transform 1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1649977179
transform 1 0 13892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_5
timestamp 1649977179
transform 1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1649977179
transform 1 0 18032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_188
timestamp 1649977179
transform 1 0 18400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_218
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1649977179
transform 1 0 13248 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_136
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_148
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1649977179
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_17
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_21
timestamp 1649977179
transform 1 0 3036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_39
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_43
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_60
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_72
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1649977179
transform 1 0 12328 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_182
timestamp 1649977179
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_61
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_76
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1649977179
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1649977179
transform 1 0 19872 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_208
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_42
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1649977179
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_110
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_146
timestamp 1649977179
transform 1 0 14536 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_182
timestamp 1649977179
transform 1 0 17848 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1649977179
transform 1 0 2024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_18
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_44
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_117
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_195
timestamp 1649977179
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_60
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_213
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1649977179
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_20
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1649977179
transform 1 0 3496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_80
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_133
timestamp 1649977179
transform 1 0 13340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1649977179
transform 1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1649977179
transform 1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_34
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1649977179
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_120
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_132
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_211
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_217
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_29
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1649977179
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_173
timestamp 1649977179
transform 1 0 17020 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1649977179
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1649977179
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_119
timestamp 1649977179
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1649977179
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1649977179
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_214
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1649977179
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_48
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_68
timestamp 1649977179
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1649977179
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_128
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_186
timestamp 1649977179
transform 1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_190
timestamp 1649977179
transform 1 0 18584 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_198
timestamp 1649977179
transform 1 0 19320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1649977179
transform 1 0 1656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_47
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1649977179
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_107
timestamp 1649977179
transform 1 0 10948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1649977179
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1649977179
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1649977179
transform 1 0 16744 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1649977179
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1649977179
transform 1 0 17480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_188
timestamp 1649977179
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_6
timestamp 1649977179
transform 1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_61
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_68
timestamp 1649977179
transform 1 0 7360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1649977179
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_100
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_104
timestamp 1649977179
transform 1 0 10672 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1649977179
transform 1 0 12420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_144
timestamp 1649977179
transform 1 0 14352 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_163
timestamp 1649977179
transform 1 0 16100 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_171
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_177
timestamp 1649977179
transform 1 0 17388 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_190
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1649977179
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_218
timestamp 1649977179
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1649977179
transform 1 0 21528 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1649977179
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_44
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1649977179
transform 1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_67
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1649977179
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_92
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_96
timestamp 1649977179
transform 1 0 9936 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_155
timestamp 1649977179
transform 1 0 15364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1649977179
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1649977179
transform 1 0 20056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1649977179
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_6
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1649977179
transform 1 0 2208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_22
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1649977179
transform 1 0 5520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_79
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1649977179
transform 1 0 10488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1649977179
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_154
timestamp 1649977179
transform 1 0 15272 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_186
timestamp 1649977179
transform 1 0 18216 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_198
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_210
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1649977179
transform 1 0 2208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1649977179
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_47
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_59
timestamp 1649977179
transform 1 0 6532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_150
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_172
timestamp 1649977179
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_217
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_12
timestamp 1649977179
transform 1 0 2208 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_16
timestamp 1649977179
transform 1 0 2576 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_76
timestamp 1649977179
transform 1 0 8096 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_124
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1649977179
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_147
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_186
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_190
timestamp 1649977179
transform 1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_206
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_212
timestamp 1649977179
transform 1 0 20608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1649977179
transform -1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform 1 0 16744 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform 1 0 12512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform -1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform 1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1649977179
transform -1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1649977179
transform -1 0 2024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1649977179
transform -1 0 2944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1649977179
transform -1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1649977179
transform -1 0 5612 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1649977179
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1649977179
transform -1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1649977179
transform -1 0 2668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform -1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform -1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform -1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform -1 0 2760 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform -1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform -1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform 1 0 20792 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform 1 0 13616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1649977179
transform -1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1649977179
transform -1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1649977179
transform -1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1649977179
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11040 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12052 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13340 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10580 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12144 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10212 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16652 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20424 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 18676 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12052 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13708 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11776 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15456 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13892 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21344 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21252 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18584 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16928 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 19872 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17572 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6440 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5980 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8280 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8556 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8004 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7912 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7360 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12420 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13432 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10672 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11684 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4876 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2760 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2760 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 1564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1840 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4692 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3588 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3864 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3680 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21252 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 19964 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 9384 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 16192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 18768 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 20332 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 12696 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform -1 0 18584 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 21068 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 17940 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21344 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6992 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12420 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14628 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14536 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15088 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
<< labels >>
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 0 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 134 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 135 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 136 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 137 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 138 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 139 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 140 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 141 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 left_top_grid_pin_1_
port 142 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 143 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 144 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 145 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 146 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 147 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 148 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 149 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 150 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 151 nsew signal input
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 right_top_grid_pin_1_
port 152 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
