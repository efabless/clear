* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

.subckt sb_1__0_ SC_IN_TOP SC_OUT_TOP Test_en_N_out Test_en_S_in ccff_head ccff_tail
+ chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13]
+ chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18]
+ chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9]
+ chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
+ chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9]
+ chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13]
+ chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18]
+ chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9]
+ chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] clk_3_N_out clk_3_S_in left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk_0_N_in
+ prog_clk_3_N_out prog_clk_3_S_in right_bottom_grid_pin_11_ right_bottom_grid_pin_13_
+ right_bottom_grid_pin_15_ right_bottom_grid_pin_17_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_
+ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_42_
+ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_
+ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_ VPWR VGND
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ _062_/A VGND VGND VPWR VPWR _062_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input55_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__buf_1
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_10.mux_l2_in_1_ _031_/HI _087_/A mux_top_track_10.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input18_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_028_ VGND VGND VPWR VPWR _028_/HI _028_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 _068_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__clkbuf_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input85_A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_061_ _061_/A VGND VGND VPWR VPWR _061_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _061_/A sky130_fd_sc_hd__clkbuf_1
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__buf_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_10.mux_l2_in_0_ input34/X mux_top_track_10.mux_l1_in_0_/X mux_top_track_10.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 _069_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__clkbuf_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_3_ _029_/HI _094_/A mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input30_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l2_in_3_ _030_/HI _080_/A mux_top_track_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input78_A right_bottom_grid_pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_mem_left_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_left_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_060_ _060_/A VGND VGND VPWR VPWR _060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__buf_1
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input60_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput99 _070_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_8.mux_l2_in_2_ _084_/A input78/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input23_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ input4/X _060_/A mux_top_track_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_10.mux_l1_in_0_ _067_/A _110_/A mux_top_track_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__064__A _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input90_A top_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmux_top_track_22.mux_l1_in_1_ _038_/HI _095_/A mux_top_track_22.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_22.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input53_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__buf_1
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__072__A _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_3_N_FTB01 input74/X VGND VGND VPWR VPWR output156/A sky130_fd_sc_hd__buf_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__067__A _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ input35/X input90/X mux_top_track_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ input83/X input79/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input16_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input8_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__080__A _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input83_A right_bottom_grid_pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l1_in_0_ _075_/A input91/X mux_top_track_22.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input46_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ input88/X mux_top_track_0.mux_l1_in_0_/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ input51/X mux_right_track_8.mux_l1_in_0_/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input76_A right_bottom_grid_pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
XANTENNA_input39_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _116_/A sky130_fd_sc_hd__buf_1
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_0_ input63/X input56/X mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l1_in_0_ input86/X input84/X mux_top_track_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A left_bottom_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input51_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_6_ _092_/A _083_/A rebuffer2/A VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_6_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input14_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input6_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l2_in_3_ _047_/HI input67/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input81_A right_bottom_grid_pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input44_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_5_ input78/X input77/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _059_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l2_in_2_ input65/X input72/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input74_A prog_clk_3_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l2_in_3_ _028_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__buf_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input37_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ input76/X input75/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l2_in_1_ input70/X _071_/A mux_left_track_3.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_6.mux_l1_in_3__A1 _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input67_A left_bottom_grid_pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l1_in_3_ _052_/HI _095_/A mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_ _034_/HI _091_/A mux_top_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_3_ input83/X input82/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_2_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l2_in_0_ _062_/A mux_left_track_3.mux_l1_in_0_/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_2_ _086_/A input75/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_2_ input81/X input80/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_ _071_/A input88/X mux_top_track_16.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input42_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput90 top_left_grid_pin_48_ VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__buf_1
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_6.mux_l1_in_3_ _042_/HI _084_/A mux_top_track_6.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ rebuffer2/X VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_0_ input48/X input60/X mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input72_A left_bottom_grid_pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_1_ input80/X input52/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_1_ input79/X input50/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input35_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput91 top_left_grid_pin_49_ VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__buf_1
Xinput80 right_bottom_grid_pin_3_ VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output141_A _112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_2_ input26/X _064_/A mux_top_track_6.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR rebuffer2/A sky130_fd_sc_hd__dfxtp_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input65_A left_bottom_grid_pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput1 SC_IN_TOP VGND VGND VPWR VPWR _056_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A0 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_0_ input45/X input57/X mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ input62/X input55/X rebuffer2/A VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input28_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_059_ _059_/A VGND VGND VPWR VPWR _059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput81 right_bottom_grid_pin_5_ VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_1
Xinput70 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__buf_1
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_6.mux_l1_in_1_ input91/X input89/X mux_top_track_6.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input10_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A Test_en_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 Test_en_S_in VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _058_/A VGND VGND VPWR VPWR _058_/X sky130_fd_sc_hd__clkbuf_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput60 chany_top_in[6] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_1
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput82 right_bottom_grid_pin_7_ VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__buf_1
Xinput71 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_1
XANTENNA_input40_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_0_ input87/X _110_/A mux_top_track_6.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input88_A top_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _057_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 input35/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput3 ccff_head VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkbuf_1
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A left_bottom_grid_pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_mem_left_track_1.prog_clk clkbuf_2_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_5_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_057_ _057_/A VGND VGND VPWR VPWR _057_/X sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput50 chany_top_in[15] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_1
Xinput61 chany_top_in[7] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_1
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput83 right_bottom_grid_pin_9_ VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__buf_1
Xinput72 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__buf_1
XANTENNA_input33_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l2_in_3_ _050_/HI input68/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_3_ _051_/HI _090_/A mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_left_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input63_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_10.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_056_ _056_/A VGND VGND VPWR VPWR _056_/X sky130_fd_sc_hd__buf_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput51 chany_top_in[16] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__buf_1
Xinput62 chany_top_in[8] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__buf_1
Xinput84 top_left_grid_pin_42_ VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput73 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__buf_1
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput40 chanx_right_in[6] VGND VGND VPWR VPWR _064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__068__A _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input26_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_3_ _045_/HI input65/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_18.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_2_ input73/X input69/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_2_ _080_/A input78/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_12.mux_l1_in_1__A1 _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_12.mux_l1_in_1_ _032_/HI _088_/A mux_top_track_12.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput5 chanx_left_in[10] VGND VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input56_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput150 _102_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
Xinput52 chany_top_in[17] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__buf_1
Xinput63 chany_top_in[9] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_1
Xinput85 top_left_grid_pin_43_ VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 chanx_right_in[15] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput74 prog_clk_3_S_in VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__clkbuf_1
Xinput41 chanx_right_in[7] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__buf_1
XANTENNA__084__A _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_2_ input70/X _075_/A mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_9.mux_l2_in_1_ _074_/A _064_/A mux_left_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_1_ input76/X input83/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_20.mux_l1_in_1__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input86_A top_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_12.mux_l1_in_0_ _068_/A input86/X mux_top_track_12.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 chanx_left_in[11] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l1_in_3_ _036_/HI _082_/A mux_top_track_2.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput140 _111_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput151 _103_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_24.mux_l1_in_3_ _054_/HI _096_/A mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xclk_3_N_FTB01 input64/X VGND VGND VPWR VPWR output155/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output155_A output155/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_1_ _039_/HI _096_/A mux_top_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
Xinput31 chanx_right_in[16] VGND VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput20 chanx_left_in[6] VGND VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput53 chany_top_in[18] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_1
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput86 top_left_grid_pin_44_ VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__buf_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 chanx_right_in[8] VGND VGND VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_2
Xinput75 right_bottom_grid_pin_11_ VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__buf_1
Xinput64 clk_3_S_in VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_1_ _066_/A input52/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_0_ input53/X mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input31_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input79_A right_bottom_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l1_in_1_ input81/X input79/X mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput7 chanx_left_in[12] VGND VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput141 _112_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput152 _104_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput130 _082_/X VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_2.mux_l1_in_2_ _062_/A input37/X mux_top_track_2.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_2_ _087_/A input76/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input61_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_0_ _076_/A input84/X mux_top_track_24.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 chany_top_in[19] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__buf_1
Xinput87 top_left_grid_pin_45_ VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__buf_1
Xinput32 chanx_right_in[17] VGND VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_2
Xinput10 chanx_left_in[15] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput43 chanx_right_in[9] VGND VGND VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_2
Xinput76 right_bottom_grid_pin_13_ VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__buf_1
Xinput65 left_bottom_grid_pin_11_ VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__buf_1
Xinput21 chanx_left_in[7] VGND VGND VPWR VPWR _114_/A sky130_fd_sc_hd__buf_1
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ input45/X input57/X mux_left_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output92_A _056_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input24_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l1_in_0_ input46/X input58/X mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l1_in_0_ input48/X input60/X mux_right_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input91_A top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput8 chanx_left_in[13] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput120 _091_/X VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput142 _113_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput153 _105_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput131 _083_/X VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_2.mux_l1_in_1_ input91/X input89/X mux_top_track_2.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_1_ input81/X input53/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input54_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
Xinput55 chany_top_in[1] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_1
Xinput44 chany_top_in[0] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__buf_1
Xinput88 top_left_grid_pin_46_ VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__buf_1
Xinput33 chanx_right_in[18] VGND VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[16] VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput66 left_bottom_grid_pin_13_ VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__buf_1
Xinput77 right_bottom_grid_pin_15_ VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__buf_1
Xinput22 chanx_left_in[8] VGND VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_6_ input68/X input67/X rebuffer1/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input17_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_6.mux_l1_in_2__A1 _064_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input84_A top_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 chanx_left_in[14] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput121 _092_/X VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput143 _114_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_2.mux_l1_in_0_ input87/X _110_/A mux_top_track_2.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput132 _084_/X VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput110 _062_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__clkbuf_2
Xmux_right_track_24.mux_l1_in_0_ input46/X input58/X mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput154 _106_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input47_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput45 chany_top_in[10] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_1
Xinput56 chany_top_in[2] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_1
Xinput89 top_left_grid_pin_47_ VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__buf_1
Xinput34 chanx_right_in[19] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[17] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xinput23 chanx_left_in[9] VGND VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_2
Xinput67 left_bottom_grid_pin_15_ VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__buf_1
Xinput78 right_bottom_grid_pin_17_ VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__buf_1
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_5.mux_l1_in_5_ input66/X input65/X rebuffer1/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_18.mux_l1_in_1__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input77_A right_bottom_grid_pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ hold3/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput122 _093_/X VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__clkbuf_2
Xoutput155 output155/A VGND VGND VPWR VPWR clk_3_N_out sky130_fd_sc_hd__clkbuf_2
Xoutput100 _071_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__clkbuf_2
Xoutput144 _115_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _085_/X VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__clkbuf_2
Xoutput111 _063_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_3_ _049_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
Xinput46 chany_top_in[11] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_1
Xinput57 chany_top_in[3] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_1
Xinput13 chanx_left_in[18] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_1_0_mem_left_track_1.prog_clk clkbuf_3_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_1_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xinput79 right_bottom_grid_pin_1_ VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__buf_1
Xinput68 left_bottom_grid_pin_17_ VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__buf_1
Xinput24 chanx_right_in[0] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 chanx_right_in[1] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__buf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_4_ input73/X input72/X rebuffer1/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input22_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_mem_left_track_1.prog_clk clkbuf_3_5_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_4_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput123 _094_/X VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput156 output156/A VGND VGND VPWR VPWR prog_clk_3_N_out sky130_fd_sc_hd__clkbuf_2
Xoutput101 _072_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput145 _116_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput134 _086_/X VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput112 _064_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xinput14 chanx_left_in[19] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_right_in[10] VGND VGND VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_2
Xinput36 chanx_right_in[2] VGND VGND VPWR VPWR _060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput47 chany_top_in[12] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__buf_1
Xinput58 chany_top_in[4] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_2
Xinput69 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_1
XANTENNA_input52_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_032_ VGND VGND VPWR VPWR _032_/HI _032_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_3_ input71/X input70/X rebuffer1/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_7_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _065_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input15_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_38.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A right_bottom_grid_pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput124 _095_/X VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput146 _098_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput135 _097_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput102 _073_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__clkbuf_2
Xoutput113 _065_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput48 chany_top_in[13] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__buf_1
Xinput59 chany_top_in[5] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_1
Xinput26 chanx_right_in[11] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__buf_1
Xinput15 chanx_left_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_1
Xinput37 chanx_right_in[3] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
X_031_ VGND VGND VPWR VPWR _031_/HI _031_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input45_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_3_ _046_/HI input66/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_2_ input69/X _072_/A rebuffer1/A VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR output94/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_18.mux_l1_in_1_ _035_/HI _092_/A mux_top_track_18.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_18.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_20.mux_l1_in_1_ _037_/HI _094_/A mux_top_track_20.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_20.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_38.mux_l1_in_0__A0 input15/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input75_A right_bottom_grid_pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput125 _096_/X VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _107_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput147 _099_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput103 _074_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput114 _066_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput49 chany_top_in[14] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__buf_1
Xinput27 chanx_right_in[12] VGND VGND VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 chanx_left_in[2] VGND VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_2
Xinput38 chanx_right_in[4] VGND VGND VPWR VPWR _062_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_030_ VGND VGND VPWR VPWR _030_/HI _030_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_1_ _063_/A input54/X rebuffer1/A VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input38_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_2_ input71/X _076_/A mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_output144_A _115_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_18.mux_l1_in_0_ _072_/A input89/X mux_top_track_18.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_20.mux_l1_in_0_ _074_/A input90/X mux_top_track_20.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input20_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput137 _108_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput148 _100_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput104 _075_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput126 _078_/X VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput115 _077_/X VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__clkbuf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_right_track_16.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input68_A left_bottom_grid_pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput28 chanx_right_in[13] VGND VGND VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 chanx_left_in[3] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__buf_1
Xinput39 chanx_right_in[5] VGND VGND VPWR VPWR _063_/A sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_5.mux_l1_in_0_ input47/X input59/X rebuffer1/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_25.mux_l1_in_1_ _067_/A input51/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__060__A _060_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input50_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_12.mux_l1_in_0__A0 _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_1_ _043_/HI _086_/A mux_top_track_8.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_mem_left_track_1.prog_clk clkbuf_2_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input13_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_1_ _055_/HI mux_right_track_32.mux_l1_in_2_/X mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput138 _109_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput149 _101_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput105 _076_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput116 _087_/X VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__clkbuf_2
XANTENNA__063__A _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput127 _079_/X VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_2_ _088_/A input77/X mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput29 chanx_right_in[14] VGND VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input80_A right_bottom_grid_pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[4] VGND VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_25.mux_l1_in_0_ input63/X input56/X mux_left_track_25.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_14.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ input30/X mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__066__A _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput139 _110_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput117 _088_/X VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput128 _080_/X VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput106 _058_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__clkbuf_2
Xmux_right_track_32.mux_l1_in_1_ input82/X input54/X mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput19 chanx_left_in[5] VGND VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_10.mux_l2_in_1__A1 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A left_bottom_grid_pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_top_track_12.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input36_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l2_in_3_ _044_/HI input68/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ _066_/A input84/X mux_top_track_8.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput118 _089_/X VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput129 _081_/X VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 _059_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l1_in_0_ input47/X input59/X mux_right_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input66_A left_bottom_grid_pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _058_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input29_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_2_ input66/X input73/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput119 _090_/X VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput108 _060_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__088__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l2_in_3_ _053_/HI _091_/A mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer1 rebuffer1/A VGND VGND VPWR VPWR rebuffer1/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_14.mux_l1_in_1__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input41_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ input71/X mux_left_track_1.mux_l1_in_2_/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input89_A top_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput109 _061_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_1.mux_l1_in_2_ input69/X _070_/A mux_left_track_1.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_2_ _082_/A input77/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_1__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer2 rebuffer2/A VGND VGND VPWR VPWR rebuffer2/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input71_A left_bottom_grid_pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_14.mux_l1_in_1_ _033_/HI _090_/A mux_top_track_14.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_14.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_left_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_38.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_38.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input34_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ _060_/A input49/X mux_left_track_1.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput92 _056_/X VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__clkbuf_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ input75/X input82/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input64_A clk_3_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_14.mux_l1_in_0_ _070_/A input87/X mux_top_track_14.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_38.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_3_ _041_/HI _083_/A mux_top_track_4.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A0 _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input27_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ output94/A VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput93 output93/A VGND VGND VPWR VPWR Test_en_N_out sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_1.mux_l1_in_0_ input61/X input44/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _048_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_left_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ input67/X input72/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_1_ input80/X input49/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_065_ _065_/A VGND VGND VPWR VPWR _065_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_2_ input41/X _063_/A mux_top_track_4.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_38.mux_l2_in_0_ _040_/HI mux_top_track_38.mux_l1_in_0_/X mux_top_track_38.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_mem_left_track_1.prog_clk clkbuf_3_1_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_0_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input87_A top_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 output94/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__clkbuf_2
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_left_track_1.prog_clk/X
+ rebuffer1/X VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_1_ _068_/A input50/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_0_ input61/X input44/X mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTest_en_N_FTB01 input2/X VGND VGND VPWR VPWR output93/A sky130_fd_sc_hd__buf_1
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_1
X_064_ _064_/A VGND VGND VPWR VPWR _064_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_mem_left_track_1.prog_clk clkbuf_3_3_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_3_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l1_in_1_ input90/X input88/X mux_top_track_4.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input32_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xoutput95 _057_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_left_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_38.mux_l1_in_0_ input15/X input24/X mux_top_track_38.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_38.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_left_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_mem_left_track_1.prog_clk clkbuf_3_7_0_mem_left_track_1.prog_clk/A VGND
+ VGND VPWR VPWR clkbuf_3_6_0_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR rebuffer1/A sky130_fd_sc_hd__dfxtp_4
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_33.mux_l1_in_0_ input62/X input55/X mux_left_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input62_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ _063_/A VGND VGND VPWR VPWR _063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ input86/X input84/X mux_top_track_4.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__buf_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input25_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_029_ VGND VGND VPWR VPWR _029_/HI _029_/LO sky130_fd_sc_hd__conb_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_left_track_1.prog_clk/X
+ mux_top_track_22.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 _067_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

