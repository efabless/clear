magic
tech sky130A
magscale 1 2
timestamp 1656942747
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 198 1980 22802 21004
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 386 0 442 800
rect 846 0 902 800
rect 1306 0 1362 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
<< obsm2 >>
rect 314 22144 606 22250
rect 774 22144 1066 22250
rect 1234 22144 1526 22250
rect 1694 22144 1986 22250
rect 2154 22144 2446 22250
rect 2614 22144 2906 22250
rect 3074 22144 3366 22250
rect 3534 22144 3826 22250
rect 3994 22144 4286 22250
rect 4454 22144 4746 22250
rect 4914 22144 5206 22250
rect 5374 22144 5666 22250
rect 5834 22144 6126 22250
rect 6294 22144 6586 22250
rect 6754 22144 7046 22250
rect 7214 22144 7506 22250
rect 7674 22144 7966 22250
rect 8134 22144 8426 22250
rect 8594 22144 8886 22250
rect 9054 22144 9346 22250
rect 9514 22144 9806 22250
rect 9974 22144 10266 22250
rect 10434 22144 10726 22250
rect 10894 22144 11186 22250
rect 11354 22144 11646 22250
rect 11814 22144 12106 22250
rect 12274 22144 12566 22250
rect 12734 22144 13026 22250
rect 13194 22144 13486 22250
rect 13654 22144 13946 22250
rect 14114 22144 14406 22250
rect 14574 22144 14866 22250
rect 15034 22144 15326 22250
rect 15494 22144 15786 22250
rect 15954 22144 16246 22250
rect 16414 22144 16706 22250
rect 16874 22144 17166 22250
rect 17334 22144 17626 22250
rect 17794 22144 18086 22250
rect 18254 22144 18546 22250
rect 18714 22144 19006 22250
rect 19174 22144 19466 22250
rect 19634 22144 19926 22250
rect 20094 22144 20386 22250
rect 20554 22144 20846 22250
rect 21014 22144 21306 22250
rect 21474 22144 21766 22250
rect 21934 22144 22226 22250
rect 22394 22144 22686 22250
rect 204 856 22796 22144
rect 204 734 330 856
rect 498 734 790 856
rect 958 734 1250 856
rect 1418 734 1710 856
rect 1878 734 2170 856
rect 2338 734 2630 856
rect 2798 734 3090 856
rect 3258 734 3550 856
rect 3718 734 4010 856
rect 4178 734 4470 856
rect 4638 734 4930 856
rect 5098 734 5390 856
rect 5558 734 5850 856
rect 6018 734 6310 856
rect 6478 734 6770 856
rect 6938 734 7230 856
rect 7398 734 7690 856
rect 7858 734 8150 856
rect 8318 734 8610 856
rect 8778 734 9070 856
rect 9238 734 9530 856
rect 9698 734 9990 856
rect 10158 734 10450 856
rect 10618 734 10910 856
rect 11078 734 11370 856
rect 11538 734 11830 856
rect 11998 734 12290 856
rect 12458 734 12750 856
rect 12918 734 13210 856
rect 13378 734 13670 856
rect 13838 734 14130 856
rect 14298 734 14590 856
rect 14758 734 15050 856
rect 15218 734 15510 856
rect 15678 734 15970 856
rect 16138 734 16430 856
rect 16598 734 16890 856
rect 17058 734 17350 856
rect 17518 734 17810 856
rect 17978 734 18270 856
rect 18438 734 18730 856
rect 18898 734 19190 856
rect 19358 734 19650 856
rect 19818 734 20110 856
rect 20278 734 20570 856
rect 20738 734 21030 856
rect 21198 734 21490 856
rect 21658 734 21950 856
rect 22118 734 22410 856
rect 22578 734 22796 856
<< metal3 >>
rect 0 20952 800 21072
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19320 800 19440
rect 0 18912 800 19032
rect 0 18504 800 18624
rect 0 18096 800 18216
rect 0 17688 800 17808
rect 0 17280 800 17400
rect 22200 17144 23000 17264
rect 0 16872 800 16992
rect 0 16464 800 16584
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15240 800 15360
rect 0 14832 800 14952
rect 0 14424 800 14544
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13200 800 13320
rect 0 12792 800 12912
rect 0 12384 800 12504
rect 0 11976 800 12096
rect 0 11568 800 11688
rect 0 11160 800 11280
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 0 9936 800 10056
rect 0 9528 800 9648
rect 0 9120 800 9240
rect 0 8712 800 8832
rect 0 8304 800 8424
rect 0 7896 800 8016
rect 0 7488 800 7608
rect 0 7080 800 7200
rect 0 6672 800 6792
rect 0 6264 800 6384
rect 0 5856 800 5976
rect 22200 5720 23000 5840
rect 0 5448 800 5568
rect 0 5040 800 5160
rect 0 4632 800 4752
rect 0 4224 800 4344
rect 0 3816 800 3936
rect 0 3408 800 3528
rect 0 3000 800 3120
rect 0 2592 800 2712
rect 0 2184 800 2304
rect 0 1776 800 1896
<< obsm3 >>
rect 880 20872 22200 21045
rect 800 20744 22200 20872
rect 880 20464 22200 20744
rect 800 20336 22200 20464
rect 880 20056 22200 20336
rect 800 19928 22200 20056
rect 880 19648 22200 19928
rect 800 19520 22200 19648
rect 880 19240 22200 19520
rect 800 19112 22200 19240
rect 880 18832 22200 19112
rect 800 18704 22200 18832
rect 880 18424 22200 18704
rect 800 18296 22200 18424
rect 880 18016 22200 18296
rect 800 17888 22200 18016
rect 880 17608 22200 17888
rect 800 17480 22200 17608
rect 880 17344 22200 17480
rect 880 17200 22120 17344
rect 800 17072 22120 17200
rect 880 17064 22120 17072
rect 880 16792 22200 17064
rect 800 16664 22200 16792
rect 880 16384 22200 16664
rect 800 16256 22200 16384
rect 880 15976 22200 16256
rect 800 15848 22200 15976
rect 880 15568 22200 15848
rect 800 15440 22200 15568
rect 880 15160 22200 15440
rect 800 15032 22200 15160
rect 880 14752 22200 15032
rect 800 14624 22200 14752
rect 880 14344 22200 14624
rect 800 14216 22200 14344
rect 880 13936 22200 14216
rect 800 13808 22200 13936
rect 880 13528 22200 13808
rect 800 13400 22200 13528
rect 880 13120 22200 13400
rect 800 12992 22200 13120
rect 880 12712 22200 12992
rect 800 12584 22200 12712
rect 880 12304 22200 12584
rect 800 12176 22200 12304
rect 880 11896 22200 12176
rect 800 11768 22200 11896
rect 880 11488 22200 11768
rect 800 11360 22200 11488
rect 880 11080 22200 11360
rect 800 10952 22200 11080
rect 880 10672 22200 10952
rect 800 10544 22200 10672
rect 880 10264 22200 10544
rect 800 10136 22200 10264
rect 880 9856 22200 10136
rect 800 9728 22200 9856
rect 880 9448 22200 9728
rect 800 9320 22200 9448
rect 880 9040 22200 9320
rect 800 8912 22200 9040
rect 880 8632 22200 8912
rect 800 8504 22200 8632
rect 880 8224 22200 8504
rect 800 8096 22200 8224
rect 880 7816 22200 8096
rect 800 7688 22200 7816
rect 880 7408 22200 7688
rect 800 7280 22200 7408
rect 880 7000 22200 7280
rect 800 6872 22200 7000
rect 880 6592 22200 6872
rect 800 6464 22200 6592
rect 880 6184 22200 6464
rect 800 6056 22200 6184
rect 880 5920 22200 6056
rect 880 5776 22120 5920
rect 800 5648 22120 5776
rect 880 5640 22120 5648
rect 880 5368 22200 5640
rect 800 5240 22200 5368
rect 880 4960 22200 5240
rect 800 4832 22200 4960
rect 880 4552 22200 4832
rect 800 4424 22200 4552
rect 880 4144 22200 4424
rect 800 4016 22200 4144
rect 880 3736 22200 4016
rect 800 3608 22200 3736
rect 880 3328 22200 3608
rect 800 3200 22200 3328
rect 880 2920 22200 3200
rect 800 2792 22200 2920
rect 880 2512 22200 2792
rect 800 2384 22200 2512
rect 880 2104 22200 2384
rect 800 1976 22200 2104
rect 880 1803 22200 1976
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 2819 2483 3463 19685
rect 3943 2483 6062 19685
rect 6542 2483 8661 19685
rect 9141 2483 11260 19685
rect 11740 2483 12085 19685
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 386 0 442 800 6 bottom_left_grid_pin_42_
port 3 nsew signal input
rlabel metal2 s 846 0 902 800 6 bottom_left_grid_pin_43_
port 4 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 bottom_left_grid_pin_44_
port 5 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 bottom_left_grid_pin_45_
port 6 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_46_
port 7 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 bottom_left_grid_pin_47_
port 8 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 bottom_left_grid_pin_48_
port 9 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 bottom_left_grid_pin_49_
port 10 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 bottom_right_grid_pin_1_
port 11 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 12 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 13 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 chanx_left_in[0]
port 14 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[10]
port 15 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 chanx_left_in[11]
port 16 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 17 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 18 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[14]
port 19 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[15]
port 20 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[16]
port 21 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[17]
port 22 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 chanx_left_in[18]
port 23 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 24 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 chanx_left_in[1]
port 25 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[2]
port 26 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[3]
port 27 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[4]
port 28 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[5]
port 29 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 chanx_left_in[6]
port 30 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 chanx_left_in[7]
port 31 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[8]
port 32 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[9]
port 33 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 34 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[10]
port 35 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 chanx_left_out[11]
port 36 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 chanx_left_out[12]
port 37 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 chanx_left_out[13]
port 38 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 chanx_left_out[14]
port 39 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[15]
port 40 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[16]
port 41 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[17]
port 42 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 chanx_left_out[18]
port 43 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 chanx_left_out[19]
port 44 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 chanx_left_out[1]
port 45 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[2]
port 46 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[3]
port 47 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 chanx_left_out[4]
port 48 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 chanx_left_out[5]
port 49 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 chanx_left_out[6]
port 50 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[7]
port 51 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[8]
port 52 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[9]
port 53 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_in[0]
port 54 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[10]
port 55 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 chany_bottom_in[11]
port 56 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 57 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[13]
port 58 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[14]
port 59 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[15]
port 60 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[16]
port 61 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[17]
port 62 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[18]
port 63 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[19]
port 64 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[1]
port 65 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[2]
port 66 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[3]
port 67 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[4]
port 68 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[5]
port 69 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[6]
port 70 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[7]
port 71 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[8]
port 72 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 chany_bottom_in[9]
port 73 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[0]
port 74 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[10]
port 75 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 chany_bottom_out[11]
port 76 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[12]
port 77 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 chany_bottom_out[13]
port 78 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 chany_bottom_out[14]
port 79 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 chany_bottom_out[15]
port 80 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[16]
port 81 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 chany_bottom_out[17]
port 82 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[18]
port 83 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 chany_bottom_out[19]
port 84 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[1]
port 85 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 chany_bottom_out[2]
port 86 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 chany_bottom_out[3]
port 87 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[4]
port 88 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 chany_bottom_out[5]
port 89 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[6]
port 90 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[7]
port 91 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[8]
port 92 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[9]
port 93 nsew signal output
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 94 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 95 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 96 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 97 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 98 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 99 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 100 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 101 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 102 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 103 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 104 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 105 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 106 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 107 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 108 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 109 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 110 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 111 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 112 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 113 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 114 nsew signal output
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 115 nsew signal output
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 116 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 117 nsew signal output
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 118 nsew signal output
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 119 nsew signal output
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 120 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 121 nsew signal output
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 122 nsew signal output
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 123 nsew signal output
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 124 nsew signal output
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 125 nsew signal output
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 126 nsew signal output
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 127 nsew signal output
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 128 nsew signal output
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 129 nsew signal output
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 130 nsew signal output
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 131 nsew signal output
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 132 nsew signal output
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 133 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 left_bottom_grid_pin_34_
port 134 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_bottom_grid_pin_35_
port 135 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 left_bottom_grid_pin_36_
port 136 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_37_
port 137 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_38_
port 138 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_39_
port 139 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 left_bottom_grid_pin_40_
port 140 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 left_bottom_grid_pin_41_
port 141 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 142 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 143 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 144 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 145 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 146 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 147 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 148 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 149 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 150 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 151 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1555434
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_2__1_/runs/sb_2__1_/results/signoff/sb_2__1_.magic.gds
string GDS_START 65026
<< end >>

