* NGSPICE file created from left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt left_tile VGND VPWR ccff_head ccff_head_0 ccff_tail ccff_tail_0 chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23]
+ chanx_right_in[24] chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28]
+ chanx_right_in[29] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21]
+ chanx_right_out[22] chanx_right_out[23] chanx_right_out[24] chanx_right_out[25]
+ chanx_right_out[26] chanx_right_out[27] chanx_right_out[28] chanx_right_out[29]
+ chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6]
+ chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2]
+ gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2]
+ gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2]
+ gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset reset right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ right_width_0_height_0_subtile_1__pin_inpad_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ right_width_0_height_0_subtile_3__pin_inpad_0_ test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_ net65 net34 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input92_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_200_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_54.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_8.mux_l1_in_0_ net73 net80 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_131_ sb_0__1_.mux_right_track_12.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input55_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_0_ net88 net73 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ sb_0__1_.mux_right_track_46.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_14.mux_l3_in_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_56.mux_l1_in_0_ net54 net105 sb_0__1_.mem_right_track_56.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_ net57 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chanx_right_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_1_ net220 net39 sb_0__1_.mem_right_track_14.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_ net71 net40 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input85_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__140__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_12.mux_l3_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_6.mux_l1_in_3_ net255 net59 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_130_ sb_0__1_.mux_right_track_14.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_52.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input48_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input102_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ sb_0__1_.mux_right_track_48.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_12.mux_l2_in_1_ net247 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0 net76 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_6.mux_l3_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_44.mux_l2_in_0__236 VGND VGND VPWR VPWR net236 sb_0__1_.mux_right_track_44.mux_l2_in_0__236/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mux_top_track_12.mux_l1_in_2_ net56 net42 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input30_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_0_ net100 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_14.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__143__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_ net78 net47 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_36.mux_l2_in_1__232 VGND VGND VPWR VPWR net232 sb_0__1_.mux_right_track_36.mux_l2_in_1__232/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input78_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_6.mux_l2_in_1_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__138__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__259 VGND VGND VPWR VPWR net259
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__259/LO sky130_fd_sc_hd__conb_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_6.mux_l1_in_2_ net46 net26 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_189_ net47 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__151__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ sb_0__1_.mux_right_track_50.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input60_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_12.mux_l2_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__146__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_3__260 VGND VGND VPWR VPWR net260 sb_0__1_.mux_top_track_0.mux_l1_in_3__260/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_12.mux_l1_in_1_ net14 net6 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__buf_2
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input23_A chanx_right_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_ net81 net50 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_26.mux_l1_in_1__227 VGND VGND VPWR VPWR net227 sb_0__1_.mux_right_track_26.mux_l1_in_1__227/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_6.mux_l2_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__154__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_14.mux_l1_in_0_ net69 net70 sb_0__1_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1 net88 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input90_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_26.mux_l2_in_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_26.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_59_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_6.mux_l1_in_1_ net8 net20 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_188_ net46 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_10.mux_l2_in_1__218 VGND VGND VPWR VPWR net218 sb_0__1_.mux_right_track_10.mux_l2_in_1__218/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_3.mux_l3_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_70_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_26.mux_l1_in_1_ net227 net60 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_111_ sb_0__1_.mux_right_track_52.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_26.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input53_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_56.mux_l2_in_0__242 VGND VGND VPWR VPWR net242 sb_0__1_.mux_right_track_56.mux_l2_in_0__242/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_30.mux_l1_in_1__229 VGND VGND VPWR VPWR net229 sb_0__1_.mux_right_track_30.mux_l1_in_1__229/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1_ net211 right_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_40.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_12.mux_l1_in_0_ net18 net107 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput101 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net101 sky130_fd_sc_hd__buf_2
XANTENNA_input16_A chanx_right_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_ sb_0__1_.mux_bottom_track_3.out
+ net53 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_36.mux_l3_in_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input8_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__170__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input83_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_1_ net251 net38 sb_0__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput202 net202 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_top_track_6.mux_l1_in_0_ net109 net107 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net111 net97 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
X_187_ sb_0__1_.mux_top_track_20.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_18.mux_l2_in_1__222 VGND VGND VPWR VPWR net222 sb_0__1_.mux_right_track_18.mux_l2_in_1__222/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_4.mux_l3_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ sb_0__1_.mux_right_track_54.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_26.mux_l1_in_0_ net106 net90 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input46_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_38.mux_l2_in_0_ net233 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_38.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input100_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_40.mux_l2_in_0_ net235 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_40.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_4.mux_l2_in_1_ net234 net47 sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__173__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_38.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net102 sky130_fd_sc_hd__buf_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__168__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_1_ net4 net16 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_top_track_4.mux_l2_in_1__252 VGND VGND VPWR VPWR net252 sb_0__1_.mux_top_track_4.mux_l2_in_1__252/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_3.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input76_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_46.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_0_ net32 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__181__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput203 net203 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_82_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_186_ net43 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__176__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input39_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_169_ net55 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_4.mux_l2_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput103 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_38.mux_l1_in_0_ net57 net104 sb_0__1_.mem_right_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__184__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_40.mux_l1_in_0_ net61 net105 sb_0__1_.mem_right_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_1_ net104 net101 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_52.mux_l2_in_0_ net240 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_52.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_right_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_0_ net92 net78 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input69_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_22.mux_l2_in_1__225 VGND VGND VPWR VPWR net225 sb_0__1_.mux_right_track_22.mux_l2_in_1__225/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.cby_0__1_.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput204 net204 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput204 net204 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3__216 VGND VGND VPWR VPWR net216 sb_0__1_.mux_bottom_track_7.mux_l1_in_3__216/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_185_ net42 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l1_in_0_ net15 net110 sb_0__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_168_ net44 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput104 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__buf_2
Xinput115 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net115 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A prog_reset_left_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_1__254 VGND VGND VPWR VPWR net254 sb_0__1_.mux_top_track_52.mux_l2_in_1__254/LO
+ sky130_fd_sc_hd__conb_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_ net258 sb_0__1_.mux_bottom_track_53.out
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_0_ net77 net83 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_38.mux_l2_in_0__233 VGND VGND VPWR VPWR net233 sb_0__1_.mux_right_track_38.mux_l2_in_0__233/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_4.mux_l2_in_1__234 VGND VGND VPWR VPWR net234 sb_0__1_.mux_right_track_4.mux_l2_in_1__234/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_44_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_29.mux_l3_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_ net64 net62 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput205 net205 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_10.mux_l3_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__257 VGND VGND VPWR VPWR net257
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__257/LO sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_right_track_52.mux_l1_in_0_ net52 net103 sb_0__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input81_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_184_ net41 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1_ net264 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_10.mux_l2_in_1_ net218 net42 sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_167_ sb_0__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net28 sb_0__1_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_right_track_0.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput105 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__buf_2
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_ net56 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_ sb_0__1_.mux_bottom_track_29.out
+ net39 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput206 net206 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XFILLER_67_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input74_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_183_ sb_0__1_.mux_top_track_28.out VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_2.mux_l3_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_top_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_10.mux_l2_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_166_ sb_0__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_22.mux_l3_in_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_22.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_1_ net10 net22 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_32.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_2.mux_l2_in_1_ net248 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0 net64 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_149_ sb_0__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput106 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_10.mux_l1_in_1_ net104 net101 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_22.mux_l2_in_1_ net225 net34 sb_0__1_.mem_right_track_22.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_1__226 VGND VGND VPWR VPWR net226 sb_0__1_.mux_right_track_24.mux_l1_in_1__226/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xleft_tile_210 VGND VGND VPWR VPWR left_tile_210/HI chanx_right_out[0] sky130_fd_sc_hd__conb_1
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_ net77 net46 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xoutput207 net207 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l3_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_23_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ net39 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input67_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_64_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_54.mux_l2_in_0__241 VGND VGND VPWR VPWR net241 sb_0__1_.mux_right_track_54.mux_l2_in_0__241/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_165_ sb_0__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l2_in_1_ net249 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_3__245 VGND VGND VPWR VPWR net245 sb_0__1_.mux_top_track_0.mux_l1_in_3__245/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_0_ net74 net69 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_30.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_2.mux_l2_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_19_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_148_ net65 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput107 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_10.mux_l1_in_0_ net72 net79 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_20.mux_l1_in_2_ net55 net41 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_22.mux_l2_in_0_ net104 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_22.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l1_in_1_ net28 net10 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input97_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_38.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input12_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_ sb_0__1_.mux_bottom_track_11.out
+ net49 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput208 net208 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input4_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_181_ net38 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_16.mux_l2_in_1__221 VGND VGND VPWR VPWR net221 sb_0__1_.mux_right_track_16.mux_l2_in_1__221/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_63_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_164_ sb_0__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_20.mux_l2_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_147_ net64 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput108 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_20.mux_l1_in_1_ net3 net5 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input42_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 chany_top_in_0[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_2.mux_l1_in_0_ net22 net108 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_4.mux_l2_in_1__249 VGND VGND VPWR VPWR net249 sb_0__1_.mux_right_track_4.mux_l2_in_1__249/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_0.mux_l3_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_22.mux_l1_in_0_ net63 net64 sb_0__1_.mem_right_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_ sb_0__1_.mux_bottom_track_5.out
+ net52 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_34.mux_l2_in_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_34.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_180_ net37 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_50.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_0.mux_l2_in_1_ net217 net51 sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input107_A top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input72_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_34.mux_l1_in_1_ net231 net55 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ net81 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_45.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_146_ net92 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput109 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__207__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_20.mux_l1_in_0_ net17 net108 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input35_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_129_ sb_0__1_.mux_right_track_16.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1__212 VGND VGND VPWR VPWR net212 sb_0__1_.mux_bottom_track_37.mux_l2_in_1__212/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput80 chany_top_in_0[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xinput91 chany_top_in_0[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_20.mux_l2_in_1__224 VGND VGND VPWR VPWR net224 sb_0__1_.mux_right_track_20.mux_l2_in_1__224/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_48.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_0.mux_l2_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_13.mux_l3_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_162_ sb_0__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input65_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_34.mux_l1_in_0_ net102 net85 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_46.mux_l2_in_0_ net237 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.mux_l2_in_1__250 VGND VGND VPWR VPWR net250 sb_0__1_.mux_top_track_28.mux_l2_in_1__250/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_right_track_0.mux_l1_in_1_ net105 net102 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_145_ sb_0__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1_ net262 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_56.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0 net71 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_128_ sb_0__1_.mux_right_track_18.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput81 chany_top_in_0[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
Xinput92 chany_top_in_0[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
Xinput70 chany_top_in_0[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_1_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ net98 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfrtp_2
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net26 sb_0__1_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input95_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_44.mux_l2_in_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input10_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A ccff_head_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_161_ sb_0__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_44.mux_l1_in_1_ net253 net37 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_6_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input58_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_24.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 ccff_head_0 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_0.mux_l1_in_0_ net99 net81 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_144_ net90 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_54.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_56.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_21_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_46.mux_l1_in_0_ net45 net100 sb_0__1_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1 net40 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_127_ sb_0__1_.mux_right_track_20.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput82 chany_top_in_0[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xinput71 chany_top_in_0[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_88_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_1_ net8 net20 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_2.mux_l2_in_1__223 VGND VGND VPWR VPWR net223 sb_0__1_.mux_right_track_2.mux_l2_in_1__223/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input40_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__144__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input88_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_ net259 net86 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__139__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ net78 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_44.mux_l1_in_0_ net31 net13 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_ net92 net61 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_22.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__152__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input105_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input70_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_20.mux_l2_in_1__249 VGND VGND VPWR VPWR net249 sb_0__1_.mux_top_track_20.mux_l2_in_1__249/LO
+ sky130_fd_sc_hd__conb_1
X_143_ net89 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__147__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_40.mux_l2_in_0__235 VGND VGND VPWR VPWR net235 sb_0__1_.mux_right_track_40.mux_l2_in_0__235/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput170 net170 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_126_ sb_0__1_.mux_right_track_22.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 chany_top_in_0[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xinput50 chany_bottom_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 chany_bottom_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 chany_top_in_0[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_0_ net86 net72 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input33_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ sb_0__1_.mux_right_track_56.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__160__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l3_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_16.mux_l3_in_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1__263 VGND VGND VPWR VPWR net263 sb_0__1_.mux_bottom_track_21.mux_l2_in_1__263/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_ net55 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__155__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1_ net212 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_1_ net221 net38 sb_0__1_.mem_right_track_16.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_52.mux_l2_in_0__240 VGND VGND VPWR VPWR net240 sb_0__1_.mux_right_track_52.mux_l2_in_0__240/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_ net69 net38 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0 net92 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ net88 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input63_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__163__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput160 net160 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ sb_0__1_.mux_right_track_24.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__158__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput73 chany_top_in_0[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput84 chany_top_in_0[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput62 chany_bottom_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput40 chany_bottom_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 chany_bottom_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XFILLER_88_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input26_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_73_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input93_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_14.mux_l2_in_1__220 VGND VGND VPWR VPWR net220 sb_0__1_.mux_right_track_14.mux_l2_in_1__220/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_37.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_0_ net101 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_16.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_ net76 net45 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1 net61 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_34.mux_l1_in_1__231 VGND VGND VPWR VPWR net231 sb_0__1_.mux_right_track_34.mux_l1_in_1__231/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_141_ sb_0__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_1_ net29 net11 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_51_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input56_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput161 net161 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
XANTENNA_input110_A top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_124_ sb_0__1_.mux_right_track_26.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__174__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput63 chany_top_in_0[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
Xinput74 chany_top_in_0[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput85 chany_top_in_0[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_right_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput52 chany_bottom_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chany_bottom_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input19_A chanx_right_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__169__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input86_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__182__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__177__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_48.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_0_ net23 net68 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_140_ net86 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input49_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_16.mux_l1_in_0_ net66 net68 sb_0__1_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput173 net173 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.mux_l2_in_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input103_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ sb_0__1_.mux_right_track_28.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 chanx_right_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 chanx_right_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_30.mux_l2_in_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_30.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput64 chany_top_in_0[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput86 chany_top_in_0[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xinput75 chany_top_in_0[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
XANTENNA__190__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput42 chany_bottom_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput53 chany_bottom_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_5.mux_l3_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA__185__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_28.mux_l1_in_1_ net228 net59 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_30.mux_l1_in_1_ net229 net58 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_90_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1_ net214 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input79_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__193__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_46.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net3 sb_0__1_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_199_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XANTENNA__188__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput174 net174 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
XFILLER_47_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input61_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__1_.mux_right_track_30.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput21 chanx_right_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 chanx_right_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chany_bottom_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput76 chany_top_in_0[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 chany_top_in_0[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput87 chany_top_in_0[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 prog_reset VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
XFILLER_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_top_track_2.mux_l2_in_1__248 VGND VGND VPWR VPWR net248 sb_0__1_.mux_top_track_2.mux_l2_in_1__248/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_right_track_6.mux_l3_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_28.mux_l1_in_0_ net99 net89 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_30.mux_l1_in_0_ net100 net88 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_90_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_right_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_6.mux_l2_in_1_ net243 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_14.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input91_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_60_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_6.mux_l1_in_2_ net46 net105 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_1_ net5 net17 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_198_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_121_ sb_0__1_.mux_right_track_32.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input54_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput88 chany_top_in_0[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput77 chany_top_in_0[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 chany_top_in_0[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_right_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_bottom_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_bottom_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
Xinput44 chany_bottom_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput99 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net99 sky130_fd_sc_hd__buf_2
XFILLER_52_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_52.mux_l3_in_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net1
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input17_A chanx_right_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_1_ net254 net35 sb_0__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input9_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_6.mux_l2_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_3__246 VGND VGND VPWR VPWR net246 sb_0__1_.mux_top_track_10.mux_l1_in_3__246/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_bottom_track_21.mux_l3_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_77_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input84_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_54.mux_l2_in_0_ net241 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_54.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_6.mux_l1_in_1_ net102 net99 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_0_ net90 net77 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_197_ sb_0__1_.mux_top_track_0.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1_ net263 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput132 net132 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
Xoutput143 net143 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput154 net154 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
XFILLER_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ sb_0__1_.mux_right_track_34.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input47_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput78 chany_top_in_0[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput67 chany_top_in_0[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput89 chany_top_in_0[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput23 chanx_right_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput56 chany_bottom_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput34 chany_bottom_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput45 chany_bottom_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input101_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net27 sb_0__1_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_34.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_0_ net30 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_29.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_6.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input77_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_6.mux_l1_in_0_ net76 net82 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ sb_0__1_.mux_top_track_2.out VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput177 net177 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_12.mux_l3_in_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_54.mux_l1_in_0_ net53 net104 sb_0__1_.mem_right_track_54.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput79 chany_top_in_0[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_top_in_0[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
X_179_ sb_0__1_.mux_top_track_36.out VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 chanx_right_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput57 chany_bottom_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chany_bottom_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3__261 VGND VGND VPWR VPWR net261 sb_0__1_.mux_bottom_track_11.mux_l1_in_3__261/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_1_ net9 net21 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_32.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_3_ net246 net58 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_12.mux_l2_in_1_ net219 net41 sb_0__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_22_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input22_A chanx_right_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_52.mux_l1_in_0_ net12 net24 sb_0__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_10.mux_l3_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_32.mux_l1_in_1__230 VGND VGND VPWR VPWR net230 sb_0__1_.mux_right_track_32.mux_l1_in_1__230/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ sb_0__1_.mux_top_track_4.out VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__258 VGND VGND VPWR VPWR net258
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__258/LO sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
Xoutput156 net156 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_top_track_10.mux_l2_in_1_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 chanx_right_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_bottom_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput69 chany_top_in_0[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
X_178_ net35 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xinput47 chany_bottom_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xinput58 chany_bottom_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_4.mux_l3_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_0_ net85 net71 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input52_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_10.mux_l1_in_2_ net43 net25 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_45.mux_l3_in_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_12.mux_l2_in_0_ net99 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_4.mux_l2_in_1_ net252 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input15_A chanx_right_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1_ net213 net30 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input7_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_6.mux_l1_in_3__255 VGND VGND VPWR VPWR net255 sb_0__1_.mux_top_track_6.mux_l1_in_3__255/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_4.mux_l1_in_2_ net60 net47 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input82_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ sb_0__1_.mux_top_track_6.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput179 net179 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_10.mux_l2_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_177_ net34 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_right_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 chanx_right_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput37 chany_bottom_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
Xinput59 chany_bottom_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
Xinput48 chany_bottom_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input45_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_10.mux_l1_in_1_ net7 net19 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1__264 VGND VGND VPWR VPWR net264 sb_0__1_.mux_bottom_track_29.mux_l2_in_1__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_4.mux_l2_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_0_ net12 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_12.mux_l1_in_0_ net71 net75 sb_0__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_24.mux_l2_in_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_24.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net2 net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mux_right_track_36.mux_l3_in_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_4.mux_l1_in_1_ net27 net9 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_82_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_50_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ net51 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input75_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1__214 VGND VGND VPWR VPWR net214 sb_0__1_.mux_bottom_track_5.mux_l2_in_1__214/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_bottom_track_1.mux_l3_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_50.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_1_ net226 net62 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput158 net158 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_36.mux_l2_in_1_ net232 net33 sb_0__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 chanx_right_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
X_176_ net62 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_right_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput38 chany_bottom_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
Xinput49 chany_bottom_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1_ net260 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input38_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_10.mux_l1_in_0_ net110 net108 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_159_ net77 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_2_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ right_width_0_height_0_subtile_0__pin_inpad_0_ sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input20_A chanx_right_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_4.mux_l1_in_0_ net21 net109 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_18.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__142__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_48.mux_l2_in_0__238 VGND VGND VPWR VPWR net238 sb_0__1_.mux_right_track_48.mux_l2_in_0__238/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_192_ sb_0__1_.mux_top_track_10.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_45.mux_l1_in_0_ net24 net67 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_2.mux_l3_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_0_ net105 net92 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xoutput159 net159 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput115 net115 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_36.mux_l2_in_0_ net44 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_175_ sb_0__1_.mux_top_track_44.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xinput17 chanx_right_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 chanx_right_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_bottom_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_0.mux_l2_in_1__217 VGND VGND VPWR VPWR net217 sb_0__1_.mux_right_track_0.mux_l2_in_1__217/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_26.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l2_in_1_ net223 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_158_ net76 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__150__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input50_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l1_in_2_ net48 net106 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_1_ net32 net15 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input98_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input13_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input5_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ sb_0__1_.mux_top_track_12.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
Xoutput116 net116 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input80_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_right_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_174_ net60 VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
Xinput29 chanx_right_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__148__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_right_track_24.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_2.mux_l2_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_157_ sb_0__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.mux_l1_in_0_ net103 net74 sb_0__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_48.mux_l2_in_0_ net238 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input43_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_50.mux_l2_in_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_50.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_2.mux_l1_in_1_ net103 net100 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_0_ net64 net81 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__156__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.out sky130_fd_sc_hd__clkbuf_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_50.mux_l1_in_1_ net239 net50 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_190_ net48 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__256 VGND VGND VPWR VPWR net256
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__256/LO sky130_fd_sc_hd__conb_1
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input108_A top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput19 chanx_right_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
X_173_ net59 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_top_track_12.mux_l2_in_1__247 VGND VGND VPWR VPWR net247 sb_0__1_.mux_top_track_12.mux_l2_in_1__247/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_8.mux_l2_in_1__244 VGND VGND VPWR VPWR net244 sb_0__1_.mux_right_track_8.mux_l2_in_1__244/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_156_ net73 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__159__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_ net256 net89 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_139_ net85 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_2.mux_l1_in_0_ net78 net84 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__172__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_48.mux_l1_in_0_ net49 net101 sb_0__1_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_ sb_0__1_.mux_bottom_track_37.out
+ net35 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_50.mux_l1_in_0_ net106 net102 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1__211 VGND VGND VPWR VPWR net211 sb_0__1_.mux_bottom_track_3.mux_l2_in_1__211/LO
+ sky130_fd_sc_hd__conb_1
Xoutput129 net129 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_23_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_172_ net58 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input66_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__180__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_155_ net72 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1__215 VGND VGND VPWR VPWR net215 sb_0__1_.mux_bottom_track_53.mux_l1_in_1__215/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input29_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_ net58 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_138_ net74 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_3_ net245 net34 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1__262 VGND VGND VPWR VPWR net262 sb_0__1_.mux_bottom_track_13.mux_l2_in_1__262/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_ net72 net41 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input96_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_40.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_0.mux_l3_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1__260 VGND VGND VPWR VPWR net260 sb_0__1_.mux_bottom_track_1.mux_l2_in_1__260/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__178__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_18.mux_l3_in_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input3_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ sb_0__1_.mux_top_track_52.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_top_track_44.mux_l1_in_1__253 VGND VGND VPWR VPWR net253 sb_0__1_.mux_top_track_44.mux_l1_in_1__253/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l3_in_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input59_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_0.mux_l2_in_1_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_154_ net71 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_50.mux_l1_in_1__239 VGND VGND VPWR VPWR net239 sb_0__1_.mux_right_track_50.mux_l1_in_1__239/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l2_in_1_ net222 net37 sb_0__1_.mem_right_track_18.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l2_in_1_ net224 net35 sb_0__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_137_ sb_0__1_.mux_right_track_0.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_2_ net51 net29 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__186__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input41_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_ sb_0__1_.mux_bottom_track_13.out
+ net48 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input89_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_170_ net56 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__189__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_0.mux_l2_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input106_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ sb_0__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input71_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l2_in_0_ net102 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_18.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_20.mux_l2_in_0_ net103 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_136_ sb_0__1_.mux_right_track_2.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
X_205_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_0.mux_l1_in_1_ net11 net23 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.out sky130_fd_sc_hd__clkbuf_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input34_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_119_ sb_0__1_.mux_right_track_36.out VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_46.mux_l2_in_0__237 VGND VGND VPWR VPWR net237 sb_0__1_.mux_right_track_46.mux_l2_in_0__237/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_66_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_28.mux_l3_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_16.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ net69 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input64_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.mux_l2_in_1_ net250 net44 sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_30.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_204_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
X_135_ sb_0__1_.mux_right_track_4.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_0_ net110 net107 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3_ net216 right_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_18.mux_l1_in_0_ net91 net67 sb_0__1_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ sb_0__1_.mux_right_track_38.out VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_20.mux_l1_in_0_ net87 net65 sb_0__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_53.mux_l2_in_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X net112 VGND VGND VPWR VPWR
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_32.mux_l2_in_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_32.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_7.mux_l3_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1_ net215 net31 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input94_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_32.mux_l1_in_1_ net230 net56 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_28.mux_l1_in_1__228 VGND VGND VPWR VPWR net228 sb_0__1_.mux_right_track_28.mux_l1_in_1__228/LO
+ sky130_fd_sc_hd__conb_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_1_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_151_ net68 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input57_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_28.mux_l2_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_203_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_134_ sb_0__1_.mux_right_track_6.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net14 sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3_ net261 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_12.mux_l2_in_1__219 VGND VGND VPWR VPWR net219 sb_0__1_.mux_right_track_12.mux_l2_in_1__219/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_28.mux_l1_in_1_ net39 net4 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_117_ sb_0__1_.mux_right_track_40.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1__213 VGND VGND VPWR VPWR net213 sb_0__1_.mux_bottom_track_45.mux_l2_in_1__213/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_8.mux_l3_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input87_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_0_ net13 net65 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_11.mux_l3_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1__275 VGND VGND VPWR VPWR net275 sb_0__1_.mux_bottom_track_1.mux_l2_in_1__275/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_32.mux_l1_in_0_ net101 net86 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_44.mux_l2_in_0_ net236 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_8.mux_l2_in_1_ net244 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_8.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_6.mux_l2_in_1__243 VGND VGND VPWR VPWR net243 sb_0__1_.mux_right_track_6.mux_l2_in_1__243/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_1_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_150_ net67 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input104_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_8.mux_l1_in_2_ net43 net106 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_133_ sb_0__1_.mux_right_track_8.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_202_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_1_ net6 net18 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net25 sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_36.mux_l2_in_1__251 VGND VGND VPWR VPWR net251 sb_0__1_.mux_top_track_36.mux_l2_in_1__251/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_top_track_28.mux_l1_in_0_ net16 net109 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ net36 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_34.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input32_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0 net81 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_8.mux_l2_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_83_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_44.mux_l1_in_0_ net40 net99 sb_0__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_8.mux_l1_in_1_ net103 net100 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_132_ sb_0__1_.mux_right_track_10.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_201_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_56.mux_l2_in_0_ net242 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_1.ccff_head VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_0_ net89 net76 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_1_ net7 net19 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_115_ sb_0__1_.mux_right_track_44.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_ net257 net88 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input25_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

