magic
tech sky130A
magscale 1 2
timestamp 1679346775
<< viali >>
rect 3249 54213 3283 54247
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10885 54213 10919 54247
rect 15485 54213 15519 54247
rect 17693 54213 17727 54247
rect 23857 54213 23891 54247
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9873 54145 9907 54179
rect 12081 54145 12115 54179
rect 14657 54145 14691 54179
rect 16313 54145 16347 54179
rect 16865 54145 16899 54179
rect 18429 54145 18463 54179
rect 19441 54145 19475 54179
rect 20269 54145 20303 54179
rect 20913 54145 20947 54179
rect 22201 54145 22235 54179
rect 22661 54145 22695 54179
rect 24777 54145 24811 54179
rect 12541 54077 12575 54111
rect 17049 54009 17083 54043
rect 20453 54009 20487 54043
rect 14841 53941 14875 53975
rect 15577 53941 15611 53975
rect 16129 53941 16163 53975
rect 17785 53941 17819 53975
rect 18521 53941 18555 53975
rect 19625 53941 19659 53975
rect 21097 53941 21131 53975
rect 22017 53941 22051 53975
rect 24593 53941 24627 53975
rect 3249 53601 3283 53635
rect 6561 53601 6595 53635
rect 8309 53601 8343 53635
rect 10517 53601 10551 53635
rect 12173 53601 12207 53635
rect 23857 53601 23891 53635
rect 2237 53533 2271 53567
rect 5457 53533 5491 53567
rect 7389 53533 7423 53567
rect 10057 53533 10091 53567
rect 11713 53533 11747 53567
rect 13737 53533 13771 53567
rect 14289 53533 14323 53567
rect 15761 53533 15795 53567
rect 16497 53533 16531 53567
rect 17417 53533 17451 53567
rect 18061 53533 18095 53567
rect 18889 53533 18923 53567
rect 19441 53533 19475 53567
rect 20545 53533 20579 53567
rect 21281 53533 21315 53567
rect 22201 53533 22235 53567
rect 22845 53533 22879 53567
rect 24777 53533 24811 53567
rect 18245 53465 18279 53499
rect 13553 53397 13587 53431
rect 14473 53397 14507 53431
rect 15945 53397 15979 53431
rect 16681 53397 16715 53431
rect 17233 53397 17267 53431
rect 18705 53397 18739 53431
rect 19625 53397 19659 53431
rect 20729 53397 20763 53431
rect 21465 53397 21499 53431
rect 22017 53397 22051 53431
rect 24593 53397 24627 53431
rect 3985 53125 4019 53159
rect 5733 53125 5767 53159
rect 14381 53125 14415 53159
rect 24869 53125 24903 53159
rect 1777 53057 1811 53091
rect 2973 53057 3007 53091
rect 4813 53057 4847 53091
rect 6837 53057 6871 53091
rect 8125 53057 8159 53091
rect 9781 53057 9815 53091
rect 11713 53057 11747 53091
rect 13553 53057 13587 53091
rect 19993 53057 20027 53091
rect 22017 53057 22051 53091
rect 22937 53057 22971 53091
rect 24133 53057 24167 53091
rect 8677 52989 8711 53023
rect 10241 52989 10275 53023
rect 12173 52989 12207 53023
rect 14565 52921 14599 52955
rect 1593 52853 1627 52887
rect 6653 52853 6687 52887
rect 13737 52853 13771 52887
rect 19809 52853 19843 52887
rect 22201 52853 22235 52887
rect 22753 52853 22787 52887
rect 11805 52649 11839 52683
rect 23765 52649 23799 52683
rect 12449 52581 12483 52615
rect 3985 52513 4019 52547
rect 4261 52513 4295 52547
rect 6101 52513 6135 52547
rect 7849 52513 7883 52547
rect 10333 52513 10367 52547
rect 2237 52445 2271 52479
rect 3249 52445 3283 52479
rect 5457 52445 5491 52479
rect 7389 52445 7423 52479
rect 9873 52445 9907 52479
rect 11989 52445 12023 52479
rect 12633 52445 12667 52479
rect 13461 52445 13495 52479
rect 23949 52445 23983 52479
rect 13277 52377 13311 52411
rect 11713 52105 11747 52139
rect 2973 51969 3007 52003
rect 4813 51969 4847 52003
rect 7113 51969 7147 52003
rect 9137 51969 9171 52003
rect 11897 51969 11931 52003
rect 25145 51969 25179 52003
rect 3525 51901 3559 51935
rect 5089 51901 5123 51935
rect 7389 51901 7423 51935
rect 9689 51901 9723 51935
rect 25237 51765 25271 51799
rect 5917 51561 5951 51595
rect 2789 51425 2823 51459
rect 4445 51425 4479 51459
rect 7021 51425 7055 51459
rect 2237 51357 2271 51391
rect 4077 51357 4111 51391
rect 6101 51357 6135 51391
rect 6745 51357 6779 51391
rect 25053 51357 25087 51391
rect 25237 51221 25271 51255
rect 6929 51017 6963 51051
rect 9873 51017 9907 51051
rect 10517 51017 10551 51051
rect 3065 50881 3099 50915
rect 6837 50881 6871 50915
rect 9781 50881 9815 50915
rect 10701 50881 10735 50915
rect 25053 50881 25087 50915
rect 1593 50813 1627 50847
rect 1869 50813 1903 50847
rect 3341 50813 3375 50847
rect 25237 50677 25271 50711
rect 6193 50473 6227 50507
rect 9413 50405 9447 50439
rect 3249 50337 3283 50371
rect 4445 50337 4479 50371
rect 2237 50269 2271 50303
rect 4077 50269 4111 50303
rect 6377 50269 6411 50303
rect 9229 50269 9263 50303
rect 25053 50269 25087 50303
rect 25237 50133 25271 50167
rect 7849 49929 7883 49963
rect 9597 49861 9631 49895
rect 1777 49793 1811 49827
rect 8033 49793 8067 49827
rect 9413 49793 9447 49827
rect 2237 49725 2271 49759
rect 2053 49249 2087 49283
rect 1593 49181 1627 49215
rect 25053 49181 25087 49215
rect 25237 49045 25271 49079
rect 11713 48841 11747 48875
rect 4261 48773 4295 48807
rect 11897 48705 11931 48739
rect 25053 48705 25087 48739
rect 3985 48637 4019 48671
rect 6009 48637 6043 48671
rect 25237 48501 25271 48535
rect 25053 48093 25087 48127
rect 1685 48025 1719 48059
rect 1869 48025 1903 48059
rect 25237 47957 25271 47991
rect 25053 47617 25087 47651
rect 25237 47413 25271 47447
rect 9137 47209 9171 47243
rect 11529 47209 11563 47243
rect 15380 47209 15414 47243
rect 15117 47073 15151 47107
rect 17877 47073 17911 47107
rect 9321 47005 9355 47039
rect 11713 47005 11747 47039
rect 17693 47005 17727 47039
rect 17785 46937 17819 46971
rect 16865 46869 16899 46903
rect 17325 46869 17359 46903
rect 7021 46665 7055 46699
rect 15393 46665 15427 46699
rect 17233 46665 17267 46699
rect 18521 46665 18555 46699
rect 17325 46597 17359 46631
rect 7205 46529 7239 46563
rect 18429 46529 18463 46563
rect 13645 46461 13679 46495
rect 13921 46461 13955 46495
rect 17417 46461 17451 46495
rect 18705 46461 18739 46495
rect 16865 46325 16899 46359
rect 18061 46325 18095 46359
rect 7757 46121 7791 46155
rect 17601 46121 17635 46155
rect 20821 46053 20855 46087
rect 16129 45985 16163 46019
rect 19901 45985 19935 46019
rect 19993 45985 20027 46019
rect 21465 45985 21499 46019
rect 1593 45917 1627 45951
rect 1869 45917 1903 45951
rect 15853 45917 15887 45951
rect 21281 45917 21315 45951
rect 25329 45917 25363 45951
rect 7665 45849 7699 45883
rect 19441 45781 19475 45815
rect 19809 45781 19843 45815
rect 21189 45781 21223 45815
rect 25145 45781 25179 45815
rect 10977 45577 11011 45611
rect 20085 45509 20119 45543
rect 20177 45509 20211 45543
rect 8585 45441 8619 45475
rect 9965 45441 9999 45475
rect 11161 45441 11195 45475
rect 11805 45441 11839 45475
rect 16865 45441 16899 45475
rect 24133 45441 24167 45475
rect 11989 45373 12023 45407
rect 13369 45373 13403 45407
rect 13645 45373 13679 45407
rect 17141 45373 17175 45407
rect 20361 45373 20395 45407
rect 24777 45373 24811 45407
rect 8401 45305 8435 45339
rect 9781 45305 9815 45339
rect 15117 45237 15151 45271
rect 18613 45237 18647 45271
rect 19717 45237 19751 45271
rect 7573 45033 7607 45067
rect 10149 45033 10183 45067
rect 16037 45033 16071 45067
rect 24593 45033 24627 45067
rect 22201 44897 22235 44931
rect 23305 44897 23339 44931
rect 23489 44897 23523 44931
rect 10701 44829 10735 44863
rect 14289 44829 14323 44863
rect 19441 44829 19475 44863
rect 23213 44829 23247 44863
rect 24777 44829 24811 44863
rect 7481 44761 7515 44795
rect 10057 44761 10091 44795
rect 10977 44761 11011 44795
rect 14565 44761 14599 44795
rect 19717 44761 19751 44795
rect 22017 44761 22051 44795
rect 22109 44761 22143 44795
rect 12449 44693 12483 44727
rect 21189 44693 21223 44727
rect 21649 44693 21683 44727
rect 22845 44693 22879 44727
rect 7297 44489 7331 44523
rect 8677 44489 8711 44523
rect 11713 44489 11747 44523
rect 14565 44489 14599 44523
rect 14657 44489 14691 44523
rect 19441 44489 19475 44523
rect 24501 44489 24535 44523
rect 7205 44353 7239 44387
rect 8033 44353 8067 44387
rect 8585 44353 8619 44387
rect 9413 44353 9447 44387
rect 12081 44353 12115 44387
rect 13001 44353 13035 44387
rect 17693 44353 17727 44387
rect 24685 44353 24719 44387
rect 25329 44353 25363 44387
rect 9689 44285 9723 44319
rect 12173 44285 12207 44319
rect 12357 44285 12391 44319
rect 14841 44285 14875 44319
rect 17969 44285 18003 44319
rect 22017 44285 22051 44319
rect 22293 44285 22327 44319
rect 7849 44217 7883 44251
rect 13185 44217 13219 44251
rect 11161 44149 11195 44183
rect 14197 44149 14231 44183
rect 23765 44149 23799 44183
rect 25145 44149 25179 44183
rect 6561 43945 6595 43979
rect 8493 43945 8527 43979
rect 9873 43945 9907 43979
rect 17601 43945 17635 43979
rect 21189 43945 21223 43979
rect 10701 43877 10735 43911
rect 16129 43809 16163 43843
rect 19717 43809 19751 43843
rect 8401 43741 8435 43775
rect 11805 43741 11839 43775
rect 15853 43741 15887 43775
rect 19441 43741 19475 43775
rect 22201 43741 22235 43775
rect 25329 43741 25363 43775
rect 6469 43673 6503 43707
rect 9781 43673 9815 43707
rect 10517 43673 10551 43707
rect 12081 43673 12115 43707
rect 22477 43673 22511 43707
rect 13553 43605 13587 43639
rect 23949 43605 23983 43639
rect 25145 43605 25179 43639
rect 5549 43401 5583 43435
rect 12265 43401 12299 43435
rect 17325 43401 17359 43435
rect 23765 43401 23799 43435
rect 5733 43265 5767 43299
rect 8585 43265 8619 43299
rect 12633 43265 12667 43299
rect 17233 43265 17267 43299
rect 24501 43265 24535 43299
rect 8861 43197 8895 43231
rect 12725 43197 12759 43231
rect 12817 43197 12851 43231
rect 17417 43197 17451 43231
rect 22017 43197 22051 43231
rect 22293 43197 22327 43231
rect 24777 43197 24811 43231
rect 10333 43061 10367 43095
rect 16865 43061 16899 43095
rect 14552 42857 14586 42891
rect 19704 42857 19738 42891
rect 4445 42721 4479 42755
rect 6561 42721 6595 42755
rect 8585 42721 8619 42755
rect 10057 42721 10091 42755
rect 12633 42721 12667 42755
rect 14289 42721 14323 42755
rect 17969 42721 18003 42755
rect 18153 42721 18187 42755
rect 19441 42721 19475 42755
rect 22293 42721 22327 42755
rect 7205 42653 7239 42687
rect 7849 42653 7883 42687
rect 9781 42653 9815 42687
rect 25329 42653 25363 42687
rect 4261 42585 4295 42619
rect 6377 42585 6411 42619
rect 8401 42585 8435 42619
rect 12357 42585 12391 42619
rect 22569 42585 22603 42619
rect 7021 42517 7055 42551
rect 7665 42517 7699 42551
rect 9413 42517 9447 42551
rect 9873 42517 9907 42551
rect 11989 42517 12023 42551
rect 12449 42517 12483 42551
rect 16037 42517 16071 42551
rect 17509 42517 17543 42551
rect 17877 42517 17911 42551
rect 21189 42517 21223 42551
rect 24041 42517 24075 42551
rect 25145 42517 25179 42551
rect 3893 42313 3927 42347
rect 11713 42313 11747 42347
rect 19625 42313 19659 42347
rect 22477 42313 22511 42347
rect 12173 42245 12207 42279
rect 21281 42245 21315 42279
rect 23581 42245 23615 42279
rect 3801 42177 3835 42211
rect 12081 42177 12115 42211
rect 17877 42177 17911 42211
rect 20545 42177 20579 42211
rect 22385 42177 22419 42211
rect 23305 42177 23339 42211
rect 7849 42109 7883 42143
rect 8125 42109 8159 42143
rect 12265 42109 12299 42143
rect 13645 42109 13679 42143
rect 13921 42109 13955 42143
rect 18153 42109 18187 42143
rect 22569 42109 22603 42143
rect 9597 41973 9631 42007
rect 15393 41973 15427 42007
rect 22017 41973 22051 42007
rect 25053 41973 25087 42007
rect 4537 41769 4571 41803
rect 7849 41769 7883 41803
rect 25145 41769 25179 41803
rect 5549 41701 5583 41735
rect 8493 41633 8527 41667
rect 11345 41633 11379 41667
rect 15301 41633 15335 41667
rect 18705 41633 18739 41667
rect 19901 41633 19935 41667
rect 20085 41633 20119 41667
rect 22109 41633 22143 41667
rect 4445 41565 4479 41599
rect 17969 41565 18003 41599
rect 21925 41565 21959 41599
rect 22017 41565 22051 41599
rect 23213 41565 23247 41599
rect 23489 41565 23523 41599
rect 25329 41565 25363 41599
rect 1685 41497 1719 41531
rect 1869 41497 1903 41531
rect 5365 41497 5399 41531
rect 11621 41497 11655 41531
rect 15577 41497 15611 41531
rect 8217 41429 8251 41463
rect 8309 41429 8343 41463
rect 13093 41429 13127 41463
rect 17049 41429 17083 41463
rect 19441 41429 19475 41463
rect 19809 41429 19843 41463
rect 21557 41429 21591 41463
rect 4077 41225 4111 41259
rect 8309 41225 8343 41259
rect 11713 41225 11747 41259
rect 12173 41225 12207 41259
rect 17325 41225 17359 41259
rect 22477 41225 22511 41259
rect 13645 41157 13679 41191
rect 17233 41157 17267 41191
rect 23489 41157 23523 41191
rect 3985 41089 4019 41123
rect 12081 41089 12115 41123
rect 13369 41089 13403 41123
rect 18429 41089 18463 41123
rect 22385 41089 22419 41123
rect 23213 41089 23247 41123
rect 6561 41021 6595 41055
rect 6837 41021 6871 41055
rect 9413 41021 9447 41055
rect 9689 41021 9723 41055
rect 12357 41021 12391 41055
rect 17417 41021 17451 41055
rect 18705 41021 18739 41055
rect 22661 41021 22695 41055
rect 11161 40885 11195 40919
rect 15117 40885 15151 40919
rect 16865 40885 16899 40919
rect 20177 40885 20211 40919
rect 21465 40885 21499 40919
rect 22017 40885 22051 40919
rect 24961 40885 24995 40919
rect 2881 40681 2915 40715
rect 17325 40681 17359 40715
rect 12817 40613 12851 40647
rect 15853 40613 15887 40647
rect 13369 40545 13403 40579
rect 16405 40545 16439 40579
rect 17877 40545 17911 40579
rect 19901 40545 19935 40579
rect 19993 40545 20027 40579
rect 21097 40545 21131 40579
rect 23857 40545 23891 40579
rect 6285 40477 6319 40511
rect 13185 40477 13219 40511
rect 16313 40477 16347 40511
rect 23765 40477 23799 40511
rect 24777 40477 24811 40511
rect 2789 40409 2823 40443
rect 6561 40409 6595 40443
rect 11437 40409 11471 40443
rect 12173 40409 12207 40443
rect 19809 40409 19843 40443
rect 21373 40409 21407 40443
rect 8033 40341 8067 40375
rect 13277 40341 13311 40375
rect 16221 40341 16255 40375
rect 17693 40341 17727 40375
rect 17785 40341 17819 40375
rect 19441 40341 19475 40375
rect 22845 40341 22879 40375
rect 23305 40341 23339 40375
rect 23673 40341 23707 40375
rect 7849 40137 7883 40171
rect 20729 40137 20763 40171
rect 21097 40137 21131 40171
rect 22017 40137 22051 40171
rect 8217 40069 8251 40103
rect 9045 40069 9079 40103
rect 9781 40069 9815 40103
rect 15577 40069 15611 40103
rect 22385 40069 22419 40103
rect 8309 40001 8343 40035
rect 22477 40001 22511 40035
rect 23213 40001 23247 40035
rect 8401 39933 8435 39967
rect 12173 39933 12207 39967
rect 12449 39933 12483 39967
rect 15669 39933 15703 39967
rect 15761 39933 15795 39967
rect 21189 39933 21223 39967
rect 21373 39933 21407 39967
rect 22569 39933 22603 39967
rect 23489 39933 23523 39967
rect 24501 39933 24535 39967
rect 13921 39797 13955 39831
rect 14565 39797 14599 39831
rect 15209 39797 15243 39831
rect 24731 39797 24765 39831
rect 7665 39593 7699 39627
rect 10596 39593 10630 39627
rect 15761 39593 15795 39627
rect 19533 39593 19567 39627
rect 20729 39593 20763 39627
rect 24593 39593 24627 39627
rect 9137 39525 9171 39559
rect 8217 39457 8251 39491
rect 9689 39457 9723 39491
rect 10333 39457 10367 39491
rect 13093 39457 13127 39491
rect 13185 39457 13219 39491
rect 14841 39457 14875 39491
rect 16405 39457 16439 39491
rect 17969 39457 18003 39491
rect 20177 39457 20211 39491
rect 21281 39457 21315 39491
rect 22385 39457 22419 39491
rect 22477 39457 22511 39491
rect 25145 39457 25179 39491
rect 9505 39389 9539 39423
rect 14749 39389 14783 39423
rect 16221 39389 16255 39423
rect 17877 39389 17911 39423
rect 21189 39389 21223 39423
rect 24041 39389 24075 39423
rect 24961 39389 24995 39423
rect 9597 39321 9631 39355
rect 14657 39321 14691 39355
rect 17785 39321 17819 39355
rect 21097 39321 21131 39355
rect 8033 39253 8067 39287
rect 8125 39253 8159 39287
rect 12081 39253 12115 39287
rect 12633 39253 12667 39287
rect 13001 39253 13035 39287
rect 14289 39253 14323 39287
rect 16129 39253 16163 39287
rect 17417 39253 17451 39287
rect 19901 39253 19935 39287
rect 19993 39253 20027 39287
rect 21925 39253 21959 39287
rect 22293 39253 22327 39287
rect 23857 39253 23891 39287
rect 25053 39253 25087 39287
rect 9689 39049 9723 39083
rect 11805 39049 11839 39083
rect 14013 39049 14047 39083
rect 15945 39049 15979 39083
rect 20361 39049 20395 39083
rect 22477 39049 22511 39083
rect 25145 39049 25179 39083
rect 10149 38981 10183 39015
rect 17969 38981 18003 39015
rect 1777 38913 1811 38947
rect 10057 38913 10091 38947
rect 12173 38913 12207 38947
rect 13185 38913 13219 38947
rect 15853 38913 15887 38947
rect 20269 38913 20303 38947
rect 22385 38913 22419 38947
rect 10241 38845 10275 38879
rect 12265 38845 12299 38879
rect 12357 38845 12391 38879
rect 14105 38845 14139 38879
rect 14289 38845 14323 38879
rect 16037 38845 16071 38879
rect 17693 38845 17727 38879
rect 20453 38845 20487 38879
rect 22569 38845 22603 38879
rect 23397 38845 23431 38879
rect 23673 38845 23707 38879
rect 13645 38777 13679 38811
rect 19441 38777 19475 38811
rect 1593 38709 1627 38743
rect 8677 38709 8711 38743
rect 11069 38709 11103 38743
rect 15485 38709 15519 38743
rect 19901 38709 19935 38743
rect 22017 38709 22051 38743
rect 6561 38505 6595 38539
rect 7849 38505 7883 38539
rect 9505 38505 9539 38539
rect 10701 38505 10735 38539
rect 16773 38505 16807 38539
rect 20637 38505 20671 38539
rect 11989 38437 12023 38471
rect 21833 38437 21867 38471
rect 4813 38369 4847 38403
rect 8493 38369 8527 38403
rect 10057 38369 10091 38403
rect 11161 38369 11195 38403
rect 11345 38369 11379 38403
rect 12449 38369 12483 38403
rect 12541 38369 12575 38403
rect 14841 38369 14875 38403
rect 14933 38369 14967 38403
rect 16313 38369 16347 38403
rect 17233 38369 17267 38403
rect 17325 38369 17359 38403
rect 19901 38369 19935 38403
rect 20085 38369 20119 38403
rect 21281 38369 21315 38403
rect 22477 38369 22511 38403
rect 23581 38369 23615 38403
rect 8217 38301 8251 38335
rect 23489 38301 23523 38335
rect 25329 38301 25363 38335
rect 5089 38233 5123 38267
rect 9965 38233 9999 38267
rect 14749 38233 14783 38267
rect 19809 38233 19843 38267
rect 21005 38233 21039 38267
rect 23397 38233 23431 38267
rect 8309 38165 8343 38199
rect 9873 38165 9907 38199
rect 11069 38165 11103 38199
rect 12357 38165 12391 38199
rect 14381 38165 14415 38199
rect 15669 38165 15703 38199
rect 15761 38165 15795 38199
rect 16129 38165 16163 38199
rect 16221 38165 16255 38199
rect 17141 38165 17175 38199
rect 19441 38165 19475 38199
rect 21097 38165 21131 38199
rect 22201 38165 22235 38199
rect 22293 38165 22327 38199
rect 23029 38165 23063 38199
rect 25145 38165 25179 38199
rect 6009 37961 6043 37995
rect 10517 37961 10551 37995
rect 12909 37961 12943 37995
rect 18797 37961 18831 37995
rect 20545 37961 20579 37995
rect 25329 37961 25363 37995
rect 13369 37893 13403 37927
rect 15393 37893 15427 37927
rect 17325 37893 17359 37927
rect 22017 37893 22051 37927
rect 23857 37893 23891 37927
rect 7573 37825 7607 37859
rect 11897 37825 11931 37859
rect 13277 37825 13311 37859
rect 14289 37825 14323 37859
rect 15301 37825 15335 37859
rect 16313 37825 16347 37859
rect 4261 37757 4295 37791
rect 4537 37757 4571 37791
rect 7849 37757 7883 37791
rect 9597 37757 9631 37791
rect 10609 37757 10643 37791
rect 10701 37757 10735 37791
rect 13553 37757 13587 37791
rect 15485 37757 15519 37791
rect 17049 37757 17083 37791
rect 20637 37757 20671 37791
rect 20729 37757 20763 37791
rect 22753 37757 22787 37791
rect 23581 37757 23615 37791
rect 10149 37689 10183 37723
rect 14933 37621 14967 37655
rect 19625 37621 19659 37655
rect 20177 37621 20211 37655
rect 5549 37281 5583 37315
rect 8309 37281 8343 37315
rect 10333 37281 10367 37315
rect 11897 37281 11931 37315
rect 15669 37281 15703 37315
rect 17049 37281 17083 37315
rect 18613 37281 18647 37315
rect 18797 37281 18831 37315
rect 21649 37281 21683 37315
rect 5273 37213 5307 37247
rect 7297 37213 7331 37247
rect 10241 37213 10275 37247
rect 15393 37213 15427 37247
rect 16773 37213 16807 37247
rect 21373 37213 21407 37247
rect 23765 37213 23799 37247
rect 24777 37213 24811 37247
rect 8125 37145 8159 37179
rect 11713 37145 11747 37179
rect 18521 37145 18555 37179
rect 19441 37145 19475 37179
rect 20177 37145 20211 37179
rect 7757 37077 7791 37111
rect 8217 37077 8251 37111
rect 9781 37077 9815 37111
rect 10149 37077 10183 37111
rect 11345 37077 11379 37111
rect 11805 37077 11839 37111
rect 15025 37077 15059 37111
rect 15485 37077 15519 37111
rect 16405 37077 16439 37111
rect 16865 37077 16899 37111
rect 17601 37077 17635 37111
rect 18153 37077 18187 37111
rect 23121 37077 23155 37111
rect 23581 37077 23615 37111
rect 24593 37077 24627 37111
rect 5181 36873 5215 36907
rect 5641 36873 5675 36907
rect 9321 36873 9355 36907
rect 12909 36873 12943 36907
rect 13369 36873 13403 36907
rect 15301 36873 15335 36907
rect 18429 36873 18463 36907
rect 19717 36873 19751 36907
rect 20177 36873 20211 36907
rect 23029 36805 23063 36839
rect 1777 36737 1811 36771
rect 5549 36737 5583 36771
rect 10149 36737 10183 36771
rect 13277 36737 13311 36771
rect 14841 36737 14875 36771
rect 15669 36737 15703 36771
rect 15761 36737 15795 36771
rect 20085 36737 20119 36771
rect 25329 36737 25363 36771
rect 5733 36669 5767 36703
rect 7573 36669 7607 36703
rect 7849 36669 7883 36703
rect 10241 36669 10275 36703
rect 10333 36669 10367 36703
rect 13461 36669 13495 36703
rect 15945 36669 15979 36703
rect 18521 36669 18555 36703
rect 18613 36669 18647 36703
rect 20269 36669 20303 36703
rect 22753 36669 22787 36703
rect 18061 36601 18095 36635
rect 1593 36533 1627 36567
rect 9781 36533 9815 36567
rect 11161 36533 11195 36567
rect 17049 36533 17083 36567
rect 24501 36533 24535 36567
rect 25145 36533 25179 36567
rect 7849 36329 7883 36363
rect 15945 36329 15979 36363
rect 21465 36329 21499 36363
rect 17141 36261 17175 36295
rect 19993 36261 20027 36295
rect 25145 36261 25179 36295
rect 6377 36193 6411 36227
rect 9873 36193 9907 36227
rect 13001 36193 13035 36227
rect 16405 36193 16439 36227
rect 16589 36193 16623 36227
rect 17693 36193 17727 36227
rect 20637 36193 20671 36227
rect 22017 36193 22051 36227
rect 23765 36193 23799 36227
rect 23949 36193 23983 36227
rect 6101 36125 6135 36159
rect 9137 36125 9171 36159
rect 11069 36125 11103 36159
rect 12909 36125 12943 36159
rect 15393 36125 15427 36159
rect 16313 36125 16347 36159
rect 17509 36125 17543 36159
rect 25329 36125 25363 36159
rect 11805 36057 11839 36091
rect 17601 36057 17635 36091
rect 20361 36057 20395 36091
rect 21925 36057 21959 36091
rect 12449 35989 12483 36023
rect 12817 35989 12851 36023
rect 20453 35989 20487 36023
rect 21833 35989 21867 36023
rect 23305 35989 23339 36023
rect 23673 35989 23707 36023
rect 6009 35785 6043 35819
rect 11161 35785 11195 35819
rect 13553 35785 13587 35819
rect 14473 35785 14507 35819
rect 15209 35785 15243 35819
rect 16865 35785 16899 35819
rect 14381 35717 14415 35751
rect 18889 35717 18923 35751
rect 23489 35717 23523 35751
rect 15577 35649 15611 35683
rect 17233 35649 17267 35683
rect 18613 35649 18647 35683
rect 22385 35649 22419 35683
rect 22477 35649 22511 35683
rect 4261 35581 4295 35615
rect 4537 35581 4571 35615
rect 9413 35581 9447 35615
rect 9689 35581 9723 35615
rect 11805 35581 11839 35615
rect 12081 35581 12115 35615
rect 14657 35581 14691 35615
rect 15669 35581 15703 35615
rect 15853 35581 15887 35615
rect 17325 35581 17359 35615
rect 17417 35581 17451 35615
rect 22569 35581 22603 35615
rect 23213 35581 23247 35615
rect 14013 35445 14047 35479
rect 20361 35445 20395 35479
rect 22017 35445 22051 35479
rect 24961 35445 24995 35479
rect 7665 35241 7699 35275
rect 9597 35241 9631 35275
rect 14841 35241 14875 35275
rect 22845 35241 22879 35275
rect 18153 35173 18187 35207
rect 25145 35173 25179 35207
rect 5549 35105 5583 35139
rect 8217 35105 8251 35139
rect 10149 35105 10183 35139
rect 12265 35105 12299 35139
rect 15301 35105 15335 35139
rect 15485 35105 15519 35139
rect 18705 35105 18739 35139
rect 20545 35105 20579 35139
rect 23397 35105 23431 35139
rect 5273 35037 5307 35071
rect 9965 35037 9999 35071
rect 11989 35037 12023 35071
rect 15209 35037 15243 35071
rect 18613 35037 18647 35071
rect 20361 35037 20395 35071
rect 25329 35037 25363 35071
rect 20453 34969 20487 35003
rect 23305 34969 23339 35003
rect 7021 34901 7055 34935
rect 8033 34901 8067 34935
rect 8125 34901 8159 34935
rect 10057 34901 10091 34935
rect 13737 34901 13771 34935
rect 18521 34901 18555 34935
rect 19993 34901 20027 34935
rect 23213 34901 23247 34935
rect 1593 34697 1627 34731
rect 5273 34697 5307 34731
rect 9045 34697 9079 34731
rect 9505 34697 9539 34731
rect 14105 34697 14139 34731
rect 14473 34697 14507 34731
rect 22017 34697 22051 34731
rect 22385 34697 22419 34731
rect 25145 34697 25179 34731
rect 7021 34629 7055 34663
rect 14565 34629 14599 34663
rect 22477 34629 22511 34663
rect 1777 34561 1811 34595
rect 3525 34561 3559 34595
rect 9413 34561 9447 34595
rect 11713 34561 11747 34595
rect 16865 34561 16899 34595
rect 19441 34561 19475 34595
rect 23397 34561 23431 34595
rect 25329 34561 25363 34595
rect 6745 34493 6779 34527
rect 9597 34493 9631 34527
rect 11989 34493 12023 34527
rect 13461 34493 13495 34527
rect 14749 34493 14783 34527
rect 17141 34493 17175 34527
rect 18613 34493 18647 34527
rect 19533 34493 19567 34527
rect 19717 34493 19751 34527
rect 22569 34493 22603 34527
rect 19073 34425 19107 34459
rect 20453 34425 20487 34459
rect 3788 34357 3822 34391
rect 8493 34357 8527 34391
rect 9137 34153 9171 34187
rect 11897 34153 11931 34187
rect 6653 34085 6687 34119
rect 5181 34017 5215 34051
rect 9689 34017 9723 34051
rect 12541 34017 12575 34051
rect 19993 34017 20027 34051
rect 21005 34017 21039 34051
rect 4905 33949 4939 33983
rect 9597 33949 9631 33983
rect 19809 33949 19843 33983
rect 20729 33949 20763 33983
rect 23857 33949 23891 33983
rect 24777 33949 24811 33983
rect 9505 33813 9539 33847
rect 12265 33813 12299 33847
rect 12357 33813 12391 33847
rect 19441 33813 19475 33847
rect 19901 33813 19935 33847
rect 22477 33813 22511 33847
rect 23673 33813 23707 33847
rect 24593 33813 24627 33847
rect 9505 33609 9539 33643
rect 9965 33609 9999 33643
rect 12265 33609 12299 33643
rect 12725 33609 12759 33643
rect 13921 33609 13955 33643
rect 15117 33609 15151 33643
rect 19533 33609 19567 33643
rect 25237 33609 25271 33643
rect 10333 33541 10367 33575
rect 13829 33541 13863 33575
rect 18613 33541 18647 33575
rect 12633 33473 12667 33507
rect 15025 33473 15059 33507
rect 18521 33473 18555 33507
rect 19901 33473 19935 33507
rect 7757 33405 7791 33439
rect 8033 33405 8067 33439
rect 10425 33405 10459 33439
rect 10517 33405 10551 33439
rect 12817 33405 12851 33439
rect 14013 33405 14047 33439
rect 15209 33405 15243 33439
rect 18705 33405 18739 33439
rect 19993 33405 20027 33439
rect 20085 33405 20119 33439
rect 23489 33405 23523 33439
rect 23765 33405 23799 33439
rect 18153 33337 18187 33371
rect 13461 33269 13495 33303
rect 14657 33269 14691 33303
rect 9137 33065 9171 33099
rect 11713 33065 11747 33099
rect 12909 33065 12943 33099
rect 18613 33065 18647 33099
rect 22109 33065 22143 33099
rect 7297 32997 7331 33031
rect 5549 32929 5583 32963
rect 9689 32929 9723 32963
rect 12265 32929 12299 32963
rect 13553 32929 13587 32963
rect 16129 32929 16163 32963
rect 16313 32929 16347 32963
rect 16865 32929 16899 32963
rect 20361 32929 20395 32963
rect 20637 32929 20671 32963
rect 23213 32929 23247 32963
rect 12081 32861 12115 32895
rect 13369 32861 13403 32895
rect 16037 32861 16071 32895
rect 19717 32861 19751 32895
rect 22937 32861 22971 32895
rect 24041 32861 24075 32895
rect 25329 32861 25363 32895
rect 5825 32793 5859 32827
rect 9505 32793 9539 32827
rect 17141 32793 17175 32827
rect 23029 32793 23063 32827
rect 9597 32725 9631 32759
rect 12173 32725 12207 32759
rect 13277 32725 13311 32759
rect 15669 32725 15703 32759
rect 19533 32725 19567 32759
rect 22569 32725 22603 32759
rect 23857 32725 23891 32759
rect 25145 32725 25179 32759
rect 17325 32521 17359 32555
rect 19441 32521 19475 32555
rect 19533 32521 19567 32555
rect 20913 32521 20947 32555
rect 23121 32521 23155 32555
rect 9413 32453 9447 32487
rect 17233 32453 17267 32487
rect 21005 32453 21039 32487
rect 1777 32385 1811 32419
rect 9137 32385 9171 32419
rect 13461 32385 13495 32419
rect 22201 32385 22235 32419
rect 23029 32385 23063 32419
rect 24041 32385 24075 32419
rect 25329 32385 25363 32419
rect 8677 32317 8711 32351
rect 14473 32317 14507 32351
rect 14749 32317 14783 32351
rect 17509 32317 17543 32351
rect 19625 32317 19659 32351
rect 21097 32317 21131 32351
rect 23213 32317 23247 32351
rect 25145 32249 25179 32283
rect 1593 32181 1627 32215
rect 7665 32181 7699 32215
rect 10885 32181 10919 32215
rect 16221 32181 16255 32215
rect 16865 32181 16899 32215
rect 19073 32181 19107 32215
rect 20545 32181 20579 32215
rect 22017 32181 22051 32215
rect 22661 32181 22695 32215
rect 23857 32181 23891 32215
rect 6929 31977 6963 32011
rect 7481 31977 7515 32011
rect 10885 31977 10919 32011
rect 12357 31977 12391 32011
rect 23857 31977 23891 32011
rect 17325 31909 17359 31943
rect 19441 31909 19475 31943
rect 20637 31909 20671 31943
rect 21833 31909 21867 31943
rect 23213 31909 23247 31943
rect 24593 31909 24627 31943
rect 5181 31841 5215 31875
rect 5457 31841 5491 31875
rect 8125 31841 8159 31875
rect 9413 31841 9447 31875
rect 12909 31841 12943 31875
rect 15117 31841 15151 31875
rect 17785 31841 17819 31875
rect 17877 31841 17911 31875
rect 21189 31841 21223 31875
rect 22477 31841 22511 31875
rect 4721 31773 4755 31807
rect 7941 31773 7975 31807
rect 9137 31773 9171 31807
rect 12817 31773 12851 31807
rect 19625 31773 19659 31807
rect 24041 31773 24075 31807
rect 24777 31773 24811 31807
rect 15393 31705 15427 31739
rect 17693 31705 17727 31739
rect 21005 31705 21039 31739
rect 21097 31705 21131 31739
rect 22201 31705 22235 31739
rect 7849 31637 7883 31671
rect 12725 31637 12759 31671
rect 16865 31637 16899 31671
rect 22293 31637 22327 31671
rect 4537 31433 4571 31467
rect 4905 31433 4939 31467
rect 7021 31433 7055 31467
rect 10149 31433 10183 31467
rect 10609 31433 10643 31467
rect 17325 31433 17359 31467
rect 4997 31365 5031 31399
rect 24869 31365 24903 31399
rect 7389 31297 7423 31331
rect 8401 31297 8435 31331
rect 10517 31297 10551 31331
rect 17693 31297 17727 31331
rect 17785 31297 17819 31331
rect 22201 31297 22235 31331
rect 23581 31297 23615 31331
rect 24685 31297 24719 31331
rect 5181 31229 5215 31263
rect 7481 31229 7515 31263
rect 7573 31229 7607 31263
rect 10701 31229 10735 31263
rect 17877 31229 17911 31263
rect 22017 31161 22051 31195
rect 23397 31093 23431 31127
rect 8401 30889 8435 30923
rect 11056 30889 11090 30923
rect 7021 30821 7055 30855
rect 13001 30821 13035 30855
rect 24869 30821 24903 30855
rect 7481 30753 7515 30787
rect 7573 30753 7607 30787
rect 10793 30753 10827 30787
rect 13553 30753 13587 30787
rect 17509 30753 17543 30787
rect 17601 30753 17635 30787
rect 22293 30753 22327 30787
rect 7389 30685 7423 30719
rect 14289 30685 14323 30719
rect 17417 30685 17451 30719
rect 14565 30617 14599 30651
rect 22569 30617 22603 30651
rect 24685 30617 24719 30651
rect 12541 30549 12575 30583
rect 13369 30549 13403 30583
rect 13461 30549 13495 30583
rect 16037 30549 16071 30583
rect 17049 30549 17083 30583
rect 24041 30549 24075 30583
rect 13093 30277 13127 30311
rect 15209 30277 15243 30311
rect 20821 30277 20855 30311
rect 20913 30277 20947 30311
rect 22385 30277 22419 30311
rect 7757 30209 7791 30243
rect 13001 30209 13035 30243
rect 17233 30209 17267 30243
rect 17325 30209 17359 30243
rect 19625 30209 19659 30243
rect 19717 30209 19751 30243
rect 23397 30209 23431 30243
rect 8033 30141 8067 30175
rect 9505 30141 9539 30175
rect 13277 30141 13311 30175
rect 15301 30141 15335 30175
rect 15393 30141 15427 30175
rect 17417 30141 17451 30175
rect 19901 30141 19935 30175
rect 21005 30141 21039 30175
rect 22477 30141 22511 30175
rect 22569 30141 22603 30175
rect 23673 30141 23707 30175
rect 12633 30073 12667 30107
rect 19257 30073 19291 30107
rect 11897 30005 11931 30039
rect 14841 30005 14875 30039
rect 16865 30005 16899 30039
rect 18705 30005 18739 30039
rect 20453 30005 20487 30039
rect 22017 30005 22051 30039
rect 25145 30005 25179 30039
rect 9137 29801 9171 29835
rect 17141 29801 17175 29835
rect 25145 29801 25179 29835
rect 11805 29733 11839 29767
rect 18061 29733 18095 29767
rect 21925 29733 21959 29767
rect 23121 29733 23155 29767
rect 2053 29665 2087 29699
rect 9781 29665 9815 29699
rect 11069 29665 11103 29699
rect 11253 29665 11287 29699
rect 12265 29665 12299 29699
rect 12357 29665 12391 29699
rect 13461 29665 13495 29699
rect 13553 29665 13587 29699
rect 17785 29665 17819 29699
rect 18613 29665 18647 29699
rect 19901 29665 19935 29699
rect 19993 29665 20027 29699
rect 21189 29665 21223 29699
rect 21373 29665 21407 29699
rect 22477 29665 22511 29699
rect 23581 29665 23615 29699
rect 23765 29665 23799 29699
rect 1777 29597 1811 29631
rect 3985 29597 4019 29631
rect 9505 29597 9539 29631
rect 10977 29597 11011 29631
rect 13369 29597 13403 29631
rect 21097 29597 21131 29631
rect 22385 29597 22419 29631
rect 25329 29597 25363 29631
rect 4169 29529 4203 29563
rect 5825 29529 5859 29563
rect 9597 29529 9631 29563
rect 18521 29529 18555 29563
rect 22293 29529 22327 29563
rect 10609 29461 10643 29495
rect 12173 29461 12207 29495
rect 13001 29461 13035 29495
rect 17509 29461 17543 29495
rect 17601 29461 17635 29495
rect 18429 29461 18463 29495
rect 19441 29461 19475 29495
rect 19809 29461 19843 29495
rect 20729 29461 20763 29495
rect 23489 29461 23523 29495
rect 9873 29257 9907 29291
rect 12265 29189 12299 29223
rect 24685 29189 24719 29223
rect 8125 29121 8159 29155
rect 12173 29121 12207 29155
rect 14565 29121 14599 29155
rect 17785 29121 17819 29155
rect 24133 29121 24167 29155
rect 12357 29053 12391 29087
rect 19533 29053 19567 29087
rect 11805 28985 11839 29019
rect 15853 28985 15887 29019
rect 23949 28985 23983 29019
rect 24869 28985 24903 29019
rect 8388 28917 8422 28951
rect 18048 28917 18082 28951
rect 22201 28917 22235 28951
rect 9137 28713 9171 28747
rect 16313 28713 16347 28747
rect 20085 28713 20119 28747
rect 21833 28713 21867 28747
rect 25145 28713 25179 28747
rect 3985 28577 4019 28611
rect 6561 28577 6595 28611
rect 9597 28577 9631 28611
rect 9689 28577 9723 28611
rect 11529 28577 11563 28611
rect 14565 28577 14599 28611
rect 14841 28577 14875 28611
rect 17509 28577 17543 28611
rect 21097 28577 21131 28611
rect 21189 28577 21223 28611
rect 22293 28577 22327 28611
rect 22477 28577 22511 28611
rect 6285 28509 6319 28543
rect 11253 28509 11287 28543
rect 17325 28509 17359 28543
rect 18337 28509 18371 28543
rect 22201 28509 22235 28543
rect 24041 28509 24075 28543
rect 25329 28509 25363 28543
rect 4169 28441 4203 28475
rect 5825 28441 5859 28475
rect 9505 28441 9539 28475
rect 8033 28373 8067 28407
rect 13001 28373 13035 28407
rect 16957 28373 16991 28407
rect 17417 28373 17451 28407
rect 20637 28373 20671 28407
rect 21005 28373 21039 28407
rect 23857 28373 23891 28407
rect 8309 28169 8343 28203
rect 10977 28169 11011 28203
rect 12357 28169 12391 28203
rect 17325 28169 17359 28203
rect 18061 28169 18095 28203
rect 22385 28169 22419 28203
rect 12449 28101 12483 28135
rect 14657 28101 14691 28135
rect 18429 28101 18463 28135
rect 18521 28101 18555 28135
rect 19809 28101 19843 28135
rect 24685 28101 24719 28135
rect 9229 28033 9263 28067
rect 14749 28033 14783 28067
rect 17233 28033 17267 28067
rect 19349 28033 19383 28067
rect 23489 28033 23523 28067
rect 24133 28033 24167 28067
rect 6561 27965 6595 27999
rect 6837 27965 6871 27999
rect 9505 27965 9539 27999
rect 12541 27965 12575 27999
rect 14841 27965 14875 27999
rect 17417 27965 17451 27999
rect 18613 27965 18647 27999
rect 19901 27965 19935 27999
rect 20085 27965 20119 27999
rect 22477 27965 22511 27999
rect 22661 27965 22695 27999
rect 11989 27897 12023 27931
rect 14289 27897 14323 27931
rect 19165 27897 19199 27931
rect 13369 27829 13403 27863
rect 16865 27829 16899 27863
rect 19441 27829 19475 27863
rect 22017 27829 22051 27863
rect 23305 27829 23339 27863
rect 23949 27829 23983 27863
rect 24777 27829 24811 27863
rect 6548 27625 6582 27659
rect 17969 27557 18003 27591
rect 24041 27557 24075 27591
rect 2053 27489 2087 27523
rect 3985 27489 4019 27523
rect 13369 27489 13403 27523
rect 14749 27489 14783 27523
rect 14933 27489 14967 27523
rect 16221 27489 16255 27523
rect 17233 27489 17267 27523
rect 17325 27489 17359 27523
rect 18429 27489 18463 27523
rect 18521 27489 18555 27523
rect 22569 27489 22603 27523
rect 1777 27421 1811 27455
rect 6285 27421 6319 27455
rect 10793 27421 10827 27455
rect 13093 27421 13127 27455
rect 17141 27421 17175 27455
rect 18337 27421 18371 27455
rect 22293 27421 22327 27455
rect 24685 27421 24719 27455
rect 4169 27353 4203 27387
rect 5825 27353 5859 27387
rect 14657 27353 14691 27387
rect 15945 27353 15979 27387
rect 24869 27353 24903 27387
rect 8033 27285 8067 27319
rect 12725 27285 12759 27319
rect 13185 27285 13219 27319
rect 14289 27285 14323 27319
rect 15577 27285 15611 27319
rect 16037 27285 16071 27319
rect 16773 27285 16807 27319
rect 2053 27081 2087 27115
rect 3479 27081 3513 27115
rect 10425 27081 10459 27115
rect 13461 27081 13495 27115
rect 17877 27081 17911 27115
rect 23949 27081 23983 27115
rect 19625 27013 19659 27047
rect 24685 27013 24719 27047
rect 2237 26945 2271 26979
rect 3408 26945 3442 26979
rect 7941 26945 7975 26979
rect 10333 26945 10367 26979
rect 11713 26945 11747 26979
rect 15025 26945 15059 26979
rect 17785 26945 17819 26979
rect 19349 26945 19383 26979
rect 8033 26877 8067 26911
rect 8125 26877 8159 26911
rect 10517 26877 10551 26911
rect 11989 26877 12023 26911
rect 15117 26877 15151 26911
rect 15209 26877 15243 26911
rect 18061 26877 18095 26911
rect 21097 26877 21131 26911
rect 22201 26877 22235 26911
rect 22477 26877 22511 26911
rect 7573 26741 7607 26775
rect 8953 26741 8987 26775
rect 9965 26741 9999 26775
rect 14657 26741 14691 26775
rect 17417 26741 17451 26775
rect 24777 26741 24811 26775
rect 8033 26537 8067 26571
rect 9321 26537 9355 26571
rect 16221 26537 16255 26571
rect 19809 26537 19843 26571
rect 23213 26537 23247 26571
rect 23857 26537 23891 26571
rect 10149 26469 10183 26503
rect 12725 26469 12759 26503
rect 3985 26401 4019 26435
rect 4905 26401 4939 26435
rect 6561 26401 6595 26435
rect 10793 26401 10827 26435
rect 13277 26401 13311 26435
rect 20361 26401 20395 26435
rect 21465 26401 21499 26435
rect 6285 26333 6319 26367
rect 10517 26333 10551 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 14473 26333 14507 26367
rect 24041 26333 24075 26367
rect 4169 26265 4203 26299
rect 10609 26265 10643 26299
rect 14749 26265 14783 26299
rect 20269 26265 20303 26299
rect 21741 26265 21775 26299
rect 24685 26265 24719 26299
rect 24869 26265 24903 26299
rect 20177 26197 20211 26231
rect 3847 25993 3881 26027
rect 7849 25993 7883 26027
rect 10425 25993 10459 26027
rect 16037 25993 16071 26027
rect 17417 25993 17451 26027
rect 19533 25993 19567 26027
rect 21281 25993 21315 26027
rect 22385 25993 22419 26027
rect 23213 25993 23247 26027
rect 10333 25925 10367 25959
rect 15117 25925 15151 25959
rect 15945 25925 15979 25959
rect 17785 25925 17819 25959
rect 24225 25925 24259 25959
rect 24961 25925 24995 25959
rect 2605 25857 2639 25891
rect 3744 25857 3778 25891
rect 19441 25857 19475 25891
rect 21465 25857 21499 25891
rect 23489 25857 23523 25891
rect 2789 25789 2823 25823
rect 7941 25789 7975 25823
rect 8033 25789 8067 25823
rect 10517 25789 10551 25823
rect 11805 25789 11839 25823
rect 12081 25789 12115 25823
rect 16221 25789 16255 25823
rect 17877 25789 17911 25823
rect 18061 25789 18095 25823
rect 19717 25789 19751 25823
rect 22477 25789 22511 25823
rect 22661 25789 22695 25823
rect 2973 25721 3007 25755
rect 7481 25721 7515 25755
rect 23673 25721 23707 25755
rect 25145 25721 25179 25755
rect 9965 25653 9999 25687
rect 13553 25653 13587 25687
rect 15577 25653 15611 25687
rect 19073 25653 19107 25687
rect 20453 25653 20487 25687
rect 22017 25653 22051 25687
rect 24317 25653 24351 25687
rect 4261 25449 4295 25483
rect 18613 25449 18647 25483
rect 12173 25381 12207 25415
rect 2053 25313 2087 25347
rect 6469 25313 6503 25347
rect 6745 25313 6779 25347
rect 12817 25313 12851 25347
rect 15577 25313 15611 25347
rect 15669 25313 15703 25347
rect 20361 25313 20395 25347
rect 20637 25313 20671 25347
rect 23029 25313 23063 25347
rect 23213 25313 23247 25347
rect 1777 25245 1811 25279
rect 3985 25245 4019 25279
rect 9321 25245 9355 25279
rect 10517 25245 10551 25279
rect 12541 25245 12575 25279
rect 13553 25245 13587 25279
rect 16865 25245 16899 25279
rect 19625 25245 19659 25279
rect 23857 25245 23891 25279
rect 24777 25245 24811 25279
rect 12633 25177 12667 25211
rect 17141 25177 17175 25211
rect 24041 25177 24075 25211
rect 4445 25109 4479 25143
rect 8217 25109 8251 25143
rect 10609 25109 10643 25143
rect 15117 25109 15151 25143
rect 15485 25109 15519 25143
rect 19441 25109 19475 25143
rect 22109 25109 22143 25143
rect 22569 25109 22603 25143
rect 22937 25109 22971 25143
rect 24593 25109 24627 25143
rect 10885 24905 10919 24939
rect 11713 24905 11747 24939
rect 12081 24905 12115 24939
rect 18337 24905 18371 24939
rect 19533 24905 19567 24939
rect 10793 24837 10827 24871
rect 2237 24769 2271 24803
rect 12173 24769 12207 24803
rect 14565 24769 14599 24803
rect 19625 24769 19659 24803
rect 22477 24769 22511 24803
rect 3065 24701 3099 24735
rect 3341 24701 3375 24735
rect 7941 24701 7975 24735
rect 8217 24701 8251 24735
rect 10977 24701 11011 24735
rect 12265 24701 12299 24735
rect 14841 24701 14875 24735
rect 16313 24701 16347 24735
rect 18429 24701 18463 24735
rect 18613 24701 18647 24735
rect 19809 24701 19843 24735
rect 22569 24701 22603 24735
rect 22753 24701 22787 24735
rect 23305 24701 23339 24735
rect 23581 24701 23615 24735
rect 2053 24633 2087 24667
rect 9689 24633 9723 24667
rect 4813 24565 4847 24599
rect 7481 24565 7515 24599
rect 10425 24565 10459 24599
rect 17969 24565 18003 24599
rect 19165 24565 19199 24599
rect 22109 24565 22143 24599
rect 25053 24565 25087 24599
rect 3157 24361 3191 24395
rect 4123 24361 4157 24395
rect 7849 24361 7883 24395
rect 14289 24361 14323 24395
rect 22201 24361 22235 24395
rect 25145 24293 25179 24327
rect 8401 24225 8435 24259
rect 9413 24225 9447 24259
rect 12173 24225 12207 24259
rect 14749 24225 14783 24259
rect 14841 24225 14875 24259
rect 15945 24225 15979 24259
rect 16129 24225 16163 24259
rect 18245 24225 18279 24259
rect 18429 24225 18463 24259
rect 19901 24225 19935 24259
rect 20085 24225 20119 24259
rect 21097 24225 21131 24259
rect 21281 24225 21315 24259
rect 2881 24157 2915 24191
rect 4020 24157 4054 24191
rect 8217 24157 8251 24191
rect 9137 24157 9171 24191
rect 11897 24157 11931 24191
rect 13737 24157 13771 24191
rect 19809 24157 19843 24191
rect 22845 24157 22879 24191
rect 25329 24157 25363 24191
rect 15853 24089 15887 24123
rect 21005 24089 21039 24123
rect 23857 24089 23891 24123
rect 3341 24021 3375 24055
rect 8309 24021 8343 24055
rect 10885 24021 10919 24055
rect 11529 24021 11563 24055
rect 11989 24021 12023 24055
rect 14657 24021 14691 24055
rect 15485 24021 15519 24055
rect 17785 24021 17819 24055
rect 18153 24021 18187 24055
rect 19441 24021 19475 24055
rect 20637 24021 20671 24055
rect 6009 23817 6043 23851
rect 8861 23817 8895 23851
rect 9689 23817 9723 23851
rect 12265 23817 12299 23851
rect 12357 23817 12391 23851
rect 13093 23817 13127 23851
rect 13461 23817 13495 23851
rect 13553 23817 13587 23851
rect 25145 23749 25179 23783
rect 2053 23681 2087 23715
rect 4261 23681 4295 23715
rect 8953 23681 8987 23715
rect 10057 23681 10091 23715
rect 11069 23681 11103 23715
rect 22293 23681 22327 23715
rect 24133 23681 24167 23715
rect 2329 23613 2363 23647
rect 9045 23613 9079 23647
rect 10149 23613 10183 23647
rect 10241 23613 10275 23647
rect 12449 23613 12483 23647
rect 13737 23613 13771 23647
rect 23305 23613 23339 23647
rect 3801 23477 3835 23511
rect 4524 23477 4558 23511
rect 8493 23477 8527 23511
rect 11897 23477 11931 23511
rect 4077 23273 4111 23307
rect 7297 23273 7331 23307
rect 15669 23205 15703 23239
rect 21005 23205 21039 23239
rect 2053 23137 2087 23171
rect 5549 23137 5583 23171
rect 10149 23137 10183 23171
rect 16313 23137 16347 23171
rect 17417 23137 17451 23171
rect 17601 23137 17635 23171
rect 21925 23137 21959 23171
rect 22017 23137 22051 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 9873 23069 9907 23103
rect 10885 23069 10919 23103
rect 16037 23069 16071 23103
rect 16129 23069 16163 23103
rect 18337 23069 18371 23103
rect 21833 23069 21867 23103
rect 22845 23069 22879 23103
rect 5825 23001 5859 23035
rect 23857 23001 23891 23035
rect 9505 22933 9539 22967
rect 9965 22933 9999 22967
rect 16957 22933 16991 22967
rect 17325 22933 17359 22967
rect 18153 22933 18187 22967
rect 21465 22933 21499 22967
rect 1961 22729 1995 22763
rect 3249 22729 3283 22763
rect 4031 22729 4065 22763
rect 12541 22729 12575 22763
rect 15117 22729 15151 22763
rect 18613 22729 18647 22763
rect 24777 22729 24811 22763
rect 7481 22661 7515 22695
rect 13645 22661 13679 22695
rect 21097 22661 21131 22695
rect 23305 22661 23339 22695
rect 2145 22593 2179 22627
rect 3928 22593 3962 22627
rect 5641 22593 5675 22627
rect 5733 22593 5767 22627
rect 15761 22593 15795 22627
rect 16865 22593 16899 22627
rect 22385 22593 22419 22627
rect 2605 22525 2639 22559
rect 2789 22525 2823 22559
rect 5917 22525 5951 22559
rect 8217 22525 8251 22559
rect 8861 22525 8895 22559
rect 9137 22525 9171 22559
rect 12633 22525 12667 22559
rect 12817 22525 12851 22559
rect 13369 22525 13403 22559
rect 19073 22525 19107 22559
rect 19349 22525 19383 22559
rect 23029 22525 23063 22559
rect 5273 22389 5307 22423
rect 10609 22389 10643 22423
rect 12173 22389 12207 22423
rect 15577 22389 15611 22423
rect 17128 22389 17162 22423
rect 22477 22389 22511 22423
rect 2697 22185 2731 22219
rect 6101 22185 6135 22219
rect 20434 22185 20468 22219
rect 14289 22117 14323 22151
rect 17417 22117 17451 22151
rect 6745 22049 6779 22083
rect 7849 22049 7883 22083
rect 11437 22049 11471 22083
rect 12449 22049 12483 22083
rect 12541 22049 12575 22083
rect 14841 22049 14875 22083
rect 15669 22049 15703 22083
rect 18613 22049 18647 22083
rect 18797 22049 18831 22083
rect 20177 22049 20211 22083
rect 2237 21981 2271 22015
rect 2881 21981 2915 22015
rect 7665 21981 7699 22015
rect 13369 21981 13403 22015
rect 14657 21981 14691 22015
rect 18521 21981 18555 22015
rect 22845 21981 22879 22015
rect 6469 21913 6503 21947
rect 10609 21913 10643 21947
rect 15945 21913 15979 21947
rect 23857 21913 23891 21947
rect 2053 21845 2087 21879
rect 6561 21845 6595 21879
rect 7297 21845 7331 21879
rect 7757 21845 7791 21879
rect 11989 21845 12023 21879
rect 12357 21845 12391 21879
rect 13185 21845 13219 21879
rect 14749 21845 14783 21879
rect 18153 21845 18187 21879
rect 21925 21845 21959 21879
rect 3157 21641 3191 21675
rect 6561 21641 6595 21675
rect 6929 21641 6963 21675
rect 7757 21641 7791 21675
rect 21373 21641 21407 21675
rect 7021 21573 7055 21607
rect 10333 21573 10367 21607
rect 14381 21573 14415 21607
rect 18153 21573 18187 21607
rect 18981 21573 19015 21607
rect 19901 21573 19935 21607
rect 22937 21573 22971 21607
rect 2513 21505 2547 21539
rect 3893 21505 3927 21539
rect 4445 21505 4479 21539
rect 8125 21505 8159 21539
rect 8217 21505 8251 21539
rect 13093 21505 13127 21539
rect 14289 21505 14323 21539
rect 15669 21505 15703 21539
rect 17509 21505 17543 21539
rect 19625 21505 19659 21539
rect 22661 21505 22695 21539
rect 2697 21437 2731 21471
rect 4905 21437 4939 21471
rect 7205 21437 7239 21471
rect 8309 21437 8343 21471
rect 10425 21437 10459 21471
rect 10609 21437 10643 21471
rect 13185 21437 13219 21471
rect 13369 21437 13403 21471
rect 14473 21437 14507 21471
rect 24685 21437 24719 21471
rect 3709 21301 3743 21335
rect 4721 21301 4755 21335
rect 9965 21301 9999 21335
rect 12725 21301 12759 21335
rect 13921 21301 13955 21335
rect 15485 21301 15519 21335
rect 3157 21097 3191 21131
rect 7665 21097 7699 21131
rect 10333 21097 10367 21131
rect 11897 21097 11931 21131
rect 13737 21097 13771 21131
rect 19441 21097 19475 21131
rect 22385 21097 22419 21131
rect 2789 20961 2823 20995
rect 3985 20961 4019 20995
rect 4261 20961 4295 20995
rect 8309 20961 8343 20995
rect 10885 20961 10919 20995
rect 12357 20961 12391 20995
rect 12541 20961 12575 20995
rect 14289 20961 14323 20995
rect 14565 20961 14599 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 20637 20961 20671 20995
rect 23397 20961 23431 20995
rect 23489 20961 23523 20995
rect 2973 20893 3007 20927
rect 10701 20893 10735 20927
rect 12265 20893 12299 20927
rect 16957 20893 16991 20927
rect 18521 20893 18555 20927
rect 19625 20893 19659 20927
rect 23305 20893 23339 20927
rect 8125 20825 8159 20859
rect 20913 20825 20947 20859
rect 5733 20757 5767 20791
rect 8033 20757 8067 20791
rect 10793 20757 10827 20791
rect 16037 20757 16071 20791
rect 18153 20757 18187 20791
rect 22937 20757 22971 20791
rect 7389 20553 7423 20587
rect 10333 20553 10367 20587
rect 12081 20553 12115 20587
rect 14749 20553 14783 20587
rect 14841 20553 14875 20587
rect 17233 20553 17267 20587
rect 17325 20553 17359 20587
rect 22385 20553 22419 20587
rect 21281 20485 21315 20519
rect 22477 20485 22511 20519
rect 23673 20485 23707 20519
rect 1777 20417 1811 20451
rect 7757 20417 7791 20451
rect 8585 20417 8619 20451
rect 15761 20417 15795 20451
rect 18797 20417 18831 20451
rect 23397 20417 23431 20451
rect 2053 20349 2087 20383
rect 7849 20349 7883 20383
rect 7941 20349 7975 20383
rect 8861 20349 8895 20383
rect 12173 20349 12207 20383
rect 12265 20349 12299 20383
rect 15025 20349 15059 20383
rect 17509 20349 17543 20383
rect 19073 20349 19107 20383
rect 22569 20349 22603 20383
rect 21465 20281 21499 20315
rect 11161 20213 11195 20247
rect 11713 20213 11747 20247
rect 14381 20213 14415 20247
rect 15577 20213 15611 20247
rect 16865 20213 16899 20247
rect 20545 20213 20579 20247
rect 22017 20213 22051 20247
rect 25145 20213 25179 20247
rect 9137 20009 9171 20043
rect 16037 20009 16071 20043
rect 4629 19873 4663 19907
rect 6101 19873 6135 19907
rect 6837 19873 6871 19907
rect 9689 19873 9723 19907
rect 11805 19873 11839 19907
rect 11989 19873 12023 19907
rect 18429 19873 18463 19907
rect 18613 19873 18647 19907
rect 21557 19873 21591 19907
rect 23857 19873 23891 19907
rect 2237 19805 2271 19839
rect 4353 19805 4387 19839
rect 6561 19805 6595 19839
rect 9505 19805 9539 19839
rect 11713 19805 11747 19839
rect 16221 19805 16255 19839
rect 17325 19805 17359 19839
rect 20729 19805 20763 19839
rect 22845 19805 22879 19839
rect 8585 19737 8619 19771
rect 17509 19737 17543 19771
rect 20085 19737 20119 19771
rect 20269 19737 20303 19771
rect 2053 19669 2087 19703
rect 9597 19669 9631 19703
rect 11345 19669 11379 19703
rect 17969 19669 18003 19703
rect 18337 19669 18371 19703
rect 4813 19465 4847 19499
rect 8125 19465 8159 19499
rect 8585 19465 8619 19499
rect 10425 19465 10459 19499
rect 13093 19465 13127 19499
rect 17877 19465 17911 19499
rect 10885 19397 10919 19431
rect 13461 19397 13495 19431
rect 17233 19397 17267 19431
rect 19441 19397 19475 19431
rect 21281 19397 21315 19431
rect 23305 19397 23339 19431
rect 4997 19329 5031 19363
rect 8493 19329 8527 19363
rect 10793 19329 10827 19363
rect 13553 19329 13587 19363
rect 18061 19329 18095 19363
rect 18705 19329 18739 19363
rect 20269 19329 20303 19363
rect 22109 19329 22143 19363
rect 24133 19329 24167 19363
rect 8769 19261 8803 19295
rect 10977 19261 11011 19295
rect 13645 19261 13679 19295
rect 24685 19261 24719 19295
rect 19625 19193 19659 19227
rect 17325 19125 17359 19159
rect 18521 19125 18555 19159
rect 3985 18921 4019 18955
rect 7205 18921 7239 18955
rect 10701 18921 10735 18955
rect 17233 18853 17267 18887
rect 21005 18853 21039 18887
rect 11345 18785 11379 18819
rect 13185 18785 13219 18819
rect 13369 18785 13403 18819
rect 17693 18785 17727 18819
rect 17877 18785 17911 18819
rect 19901 18785 19935 18819
rect 20085 18785 20119 18819
rect 21649 18785 21683 18819
rect 23949 18785 23983 18819
rect 2237 18717 2271 18751
rect 4169 18717 4203 18751
rect 5457 18717 5491 18751
rect 11069 18717 11103 18751
rect 16589 18717 16623 18751
rect 19809 18717 19843 18751
rect 21465 18717 21499 18751
rect 22201 18717 22235 18751
rect 24685 18717 24719 18751
rect 5733 18649 5767 18683
rect 17601 18649 17635 18683
rect 21373 18649 21407 18683
rect 22477 18649 22511 18683
rect 2053 18581 2087 18615
rect 11161 18581 11195 18615
rect 12725 18581 12759 18615
rect 13093 18581 13127 18615
rect 16681 18581 16715 18615
rect 19441 18581 19475 18615
rect 24777 18581 24811 18615
rect 11069 18377 11103 18411
rect 12449 18377 12483 18411
rect 12817 18377 12851 18411
rect 24501 18377 24535 18411
rect 14105 18309 14139 18343
rect 18061 18309 18095 18343
rect 23029 18309 23063 18343
rect 1777 18241 1811 18275
rect 12909 18241 12943 18275
rect 14013 18241 14047 18275
rect 19625 18241 19659 18275
rect 20269 18241 20303 18275
rect 22109 18241 22143 18275
rect 2053 18173 2087 18207
rect 6929 18173 6963 18207
rect 7205 18173 7239 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 13001 18173 13035 18207
rect 14289 18173 14323 18207
rect 18797 18173 18831 18207
rect 21281 18173 21315 18207
rect 22753 18173 22787 18207
rect 13645 18105 13679 18139
rect 8677 18037 8711 18071
rect 19441 18037 19475 18071
rect 22201 18037 22235 18071
rect 9413 17833 9447 17867
rect 17693 17833 17727 17867
rect 4813 17697 4847 17731
rect 13093 17697 13127 17731
rect 14933 17697 14967 17731
rect 15945 17697 15979 17731
rect 19717 17697 19751 17731
rect 23857 17697 23891 17731
rect 8401 17629 8435 17663
rect 9137 17629 9171 17663
rect 13001 17629 13035 17663
rect 18337 17629 18371 17663
rect 19441 17629 19475 17663
rect 22661 17629 22695 17663
rect 5089 17561 5123 17595
rect 7665 17561 7699 17595
rect 10057 17561 10091 17595
rect 10793 17561 10827 17595
rect 12909 17561 12943 17595
rect 16221 17561 16255 17595
rect 6561 17493 6595 17527
rect 9597 17493 9631 17527
rect 12541 17493 12575 17527
rect 14289 17493 14323 17527
rect 14657 17493 14691 17527
rect 14749 17493 14783 17527
rect 18429 17493 18463 17527
rect 21189 17493 21223 17527
rect 5273 17289 5307 17323
rect 5733 17289 5767 17323
rect 8677 17289 8711 17323
rect 9137 17289 9171 17323
rect 10149 17289 10183 17323
rect 12081 17289 12115 17323
rect 13645 17289 13679 17323
rect 16037 17289 16071 17323
rect 19165 17289 19199 17323
rect 21465 17289 21499 17323
rect 9045 17221 9079 17255
rect 10517 17221 10551 17255
rect 12173 17221 12207 17255
rect 14749 17221 14783 17255
rect 19993 17221 20027 17255
rect 22293 17221 22327 17255
rect 5641 17153 5675 17187
rect 7849 17153 7883 17187
rect 7941 17153 7975 17187
rect 15945 17153 15979 17187
rect 17417 17153 17451 17187
rect 19717 17153 19751 17187
rect 22017 17153 22051 17187
rect 5917 17085 5951 17119
rect 8033 17085 8067 17119
rect 9229 17085 9263 17119
rect 10609 17085 10643 17119
rect 10793 17085 10827 17119
rect 12357 17085 12391 17119
rect 13737 17085 13771 17119
rect 13921 17085 13955 17119
rect 16221 17085 16255 17119
rect 17693 17085 17727 17119
rect 13277 17017 13311 17051
rect 7481 16949 7515 16983
rect 11713 16949 11747 16983
rect 14841 16949 14875 16983
rect 15577 16949 15611 16983
rect 23765 16949 23799 16983
rect 9137 16677 9171 16711
rect 5917 16609 5951 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 10793 16609 10827 16643
rect 10977 16609 11011 16643
rect 11897 16609 11931 16643
rect 12173 16609 12207 16643
rect 22109 16609 22143 16643
rect 2513 16541 2547 16575
rect 5641 16541 5675 16575
rect 8585 16541 8619 16575
rect 9505 16541 9539 16575
rect 15945 16541 15979 16575
rect 20453 16541 20487 16575
rect 22661 16541 22695 16575
rect 23857 16541 23891 16575
rect 7665 16473 7699 16507
rect 21189 16473 21223 16507
rect 21925 16473 21959 16507
rect 2605 16405 2639 16439
rect 10333 16405 10367 16439
rect 10701 16405 10735 16439
rect 13645 16405 13679 16439
rect 15761 16405 15795 16439
rect 7021 16201 7055 16235
rect 7481 16201 7515 16235
rect 9137 16201 9171 16235
rect 9229 16201 9263 16235
rect 10793 16201 10827 16235
rect 18613 16201 18647 16235
rect 20453 16201 20487 16235
rect 21373 16201 21407 16235
rect 16129 16133 16163 16167
rect 21281 16133 21315 16167
rect 22293 16133 22327 16167
rect 1777 16065 1811 16099
rect 7389 16065 7423 16099
rect 10885 16065 10919 16099
rect 15209 16065 15243 16099
rect 16865 16065 16899 16099
rect 20361 16065 20395 16099
rect 2053 15997 2087 16031
rect 7573 15997 7607 16031
rect 9413 15997 9447 16031
rect 10977 15997 11011 16031
rect 15301 15997 15335 16031
rect 15485 15997 15519 16031
rect 17141 15997 17175 16031
rect 20545 15997 20579 16031
rect 22017 15997 22051 16031
rect 8769 15929 8803 15963
rect 16313 15929 16347 15963
rect 10425 15861 10459 15895
rect 14841 15861 14875 15895
rect 19533 15861 19567 15895
rect 19993 15861 20027 15895
rect 23765 15861 23799 15895
rect 24409 15861 24443 15895
rect 7849 15657 7883 15691
rect 11989 15657 12023 15691
rect 18153 15657 18187 15691
rect 19441 15589 19475 15623
rect 21465 15589 21499 15623
rect 6101 15521 6135 15555
rect 10517 15521 10551 15555
rect 18705 15521 18739 15555
rect 19901 15521 19935 15555
rect 20085 15521 20119 15555
rect 20821 15521 20855 15555
rect 22017 15521 22051 15555
rect 23857 15521 23891 15555
rect 10241 15453 10275 15487
rect 14381 15453 14415 15487
rect 16773 15453 16807 15487
rect 18613 15453 18647 15487
rect 22661 15453 22695 15487
rect 6377 15385 6411 15419
rect 16957 15385 16991 15419
rect 21833 15385 21867 15419
rect 14473 15317 14507 15351
rect 18521 15317 18555 15351
rect 19809 15317 19843 15351
rect 21925 15317 21959 15351
rect 7573 15113 7607 15147
rect 7941 15113 7975 15147
rect 13093 15113 13127 15147
rect 13461 15113 13495 15147
rect 19257 15113 19291 15147
rect 19625 15113 19659 15147
rect 8033 15045 8067 15079
rect 12449 15045 12483 15079
rect 13553 15045 13587 15079
rect 19717 15045 19751 15079
rect 23305 15045 23339 15079
rect 17417 14977 17451 15011
rect 18797 14977 18831 15011
rect 21005 14977 21039 15011
rect 22201 14977 22235 15011
rect 24133 14977 24167 15011
rect 8217 14909 8251 14943
rect 8769 14909 8803 14943
rect 9045 14909 9079 14943
rect 12633 14909 12667 14943
rect 13645 14909 13679 14943
rect 17509 14909 17543 14943
rect 17601 14909 17635 14943
rect 19901 14909 19935 14943
rect 24777 14909 24811 14943
rect 10517 14773 10551 14807
rect 17049 14773 17083 14807
rect 20821 14773 20855 14807
rect 9229 14569 9263 14603
rect 10682 14569 10716 14603
rect 12817 14569 12851 14603
rect 16773 14569 16807 14603
rect 6837 14433 6871 14467
rect 9873 14433 9907 14467
rect 13369 14433 13403 14467
rect 15025 14433 15059 14467
rect 10425 14365 10459 14399
rect 13185 14365 13219 14399
rect 17509 14365 17543 14399
rect 20637 14365 20671 14399
rect 23397 14365 23431 14399
rect 7113 14297 7147 14331
rect 13277 14297 13311 14331
rect 15301 14297 15335 14331
rect 18061 14297 18095 14331
rect 18245 14297 18279 14331
rect 8585 14229 8619 14263
rect 9597 14229 9631 14263
rect 9689 14229 9723 14263
rect 12173 14229 12207 14263
rect 17325 14229 17359 14263
rect 20453 14229 20487 14263
rect 23213 14229 23247 14263
rect 12725 14025 12759 14059
rect 13093 14025 13127 14059
rect 13185 14025 13219 14059
rect 13921 14025 13955 14059
rect 18613 14025 18647 14059
rect 21189 14025 21223 14059
rect 22017 14025 22051 14059
rect 9137 13957 9171 13991
rect 14289 13957 14323 13991
rect 15301 13957 15335 13991
rect 19901 13957 19935 13991
rect 21097 13957 21131 13991
rect 25145 13957 25179 13991
rect 1777 13889 1811 13923
rect 8861 13889 8895 13923
rect 10885 13889 10919 13923
rect 14381 13889 14415 13923
rect 16865 13889 16899 13923
rect 20085 13889 20119 13923
rect 22201 13889 22235 13923
rect 22845 13889 22879 13923
rect 23949 13889 23983 13923
rect 2789 13821 2823 13855
rect 13277 13821 13311 13855
rect 14565 13821 14599 13855
rect 15485 13821 15519 13855
rect 17141 13821 17175 13855
rect 21281 13821 21315 13855
rect 19257 13685 19291 13719
rect 20729 13685 20763 13719
rect 22661 13685 22695 13719
rect 18153 13481 18187 13515
rect 23305 13481 23339 13515
rect 11989 13413 12023 13447
rect 7113 13345 7147 13379
rect 12541 13345 12575 13379
rect 18613 13345 18647 13379
rect 18705 13345 18739 13379
rect 6837 13277 6871 13311
rect 12357 13277 12391 13311
rect 12449 13277 12483 13311
rect 14933 13277 14967 13311
rect 16865 13277 16899 13311
rect 18521 13277 18555 13311
rect 20913 13277 20947 13311
rect 23949 13277 23983 13311
rect 15117 13209 15151 13243
rect 19717 13209 19751 13243
rect 19901 13209 19935 13243
rect 21189 13209 21223 13243
rect 8585 13141 8619 13175
rect 22661 13141 22695 13175
rect 23765 13141 23799 13175
rect 9413 12937 9447 12971
rect 11805 12937 11839 12971
rect 16037 12937 16071 12971
rect 17233 12937 17267 12971
rect 17325 12937 17359 12971
rect 18521 12937 18555 12971
rect 21465 12937 21499 12971
rect 12265 12869 12299 12903
rect 13645 12869 13679 12903
rect 14565 12869 14599 12903
rect 19993 12869 20027 12903
rect 23305 12869 23339 12903
rect 9321 12801 9355 12835
rect 12173 12801 12207 12835
rect 14289 12801 14323 12835
rect 18429 12801 18463 12835
rect 22109 12801 22143 12835
rect 23949 12801 23983 12835
rect 9597 12733 9631 12767
rect 12357 12733 12391 12767
rect 17417 12733 17451 12767
rect 18705 12733 18739 12767
rect 19717 12733 19751 12767
rect 24777 12733 24811 12767
rect 13829 12665 13863 12699
rect 16865 12665 16899 12699
rect 8953 12597 8987 12631
rect 18061 12597 18095 12631
rect 11161 12393 11195 12427
rect 20913 12393 20947 12427
rect 16221 12325 16255 12359
rect 9689 12257 9723 12291
rect 14841 12257 14875 12291
rect 9413 12189 9447 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 16405 12189 16439 12223
rect 21097 12189 21131 12223
rect 22661 12189 22695 12223
rect 24777 12189 24811 12223
rect 13553 12121 13587 12155
rect 14749 12121 14783 12155
rect 15577 12121 15611 12155
rect 15761 12121 15795 12155
rect 17969 12121 18003 12155
rect 18153 12121 18187 12155
rect 19533 12121 19567 12155
rect 23857 12121 23891 12155
rect 13645 12053 13679 12087
rect 14289 12053 14323 12087
rect 14657 12053 14691 12087
rect 19625 12053 19659 12087
rect 24593 12053 24627 12087
rect 14381 11849 14415 11883
rect 14933 11849 14967 11883
rect 15301 11849 15335 11883
rect 18981 11849 19015 11883
rect 19625 11849 19659 11883
rect 22385 11849 22419 11883
rect 12909 11781 12943 11815
rect 16313 11713 16347 11747
rect 17233 11713 17267 11747
rect 19809 11713 19843 11747
rect 20361 11713 20395 11747
rect 22569 11713 22603 11747
rect 23397 11713 23431 11747
rect 23949 11713 23983 11747
rect 12633 11645 12667 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 17509 11645 17543 11679
rect 24685 11645 24719 11679
rect 20545 11577 20579 11611
rect 23213 11509 23247 11543
rect 13001 11305 13035 11339
rect 18153 11305 18187 11339
rect 24777 11305 24811 11339
rect 14289 11237 14323 11271
rect 19441 11237 19475 11271
rect 11253 11169 11287 11203
rect 14933 11169 14967 11203
rect 16037 11169 16071 11203
rect 19901 11169 19935 11203
rect 19993 11169 20027 11203
rect 14657 11101 14691 11135
rect 15853 11101 15887 11135
rect 18337 11101 18371 11135
rect 19809 11101 19843 11135
rect 20821 11101 20855 11135
rect 22937 11101 22971 11135
rect 24041 11101 24075 11135
rect 11529 11033 11563 11067
rect 15945 11033 15979 11067
rect 24685 11033 24719 11067
rect 14749 10965 14783 10999
rect 15485 10965 15519 10999
rect 22753 10965 22787 10999
rect 23857 10965 23891 10999
rect 19809 10761 19843 10795
rect 18337 10693 18371 10727
rect 18061 10625 18095 10659
rect 21281 10625 21315 10659
rect 23949 10625 23983 10659
rect 24777 10557 24811 10591
rect 21097 10421 21131 10455
rect 11621 10013 11655 10047
rect 16957 10013 16991 10047
rect 22845 10013 22879 10047
rect 24777 10013 24811 10047
rect 23857 9945 23891 9979
rect 11713 9877 11747 9911
rect 17049 9877 17083 9911
rect 24593 9877 24627 9911
rect 14289 9605 14323 9639
rect 6009 9537 6043 9571
rect 6929 9537 6963 9571
rect 22201 9537 22235 9571
rect 23949 9537 23983 9571
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 24777 9469 24811 9503
rect 6561 9401 6595 9435
rect 14473 9401 14507 9435
rect 22017 9333 22051 9367
rect 16129 8925 16163 8959
rect 18521 8925 18555 8959
rect 24041 8925 24075 8959
rect 24777 8925 24811 8959
rect 16313 8857 16347 8891
rect 18705 8857 18739 8891
rect 23857 8789 23891 8823
rect 24593 8789 24627 8823
rect 5917 8517 5951 8551
rect 25145 8517 25179 8551
rect 3893 8449 3927 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 4169 8381 4203 8415
rect 23305 8381 23339 8415
rect 18705 7837 18739 7871
rect 20361 7837 20395 7871
rect 22845 7837 22879 7871
rect 24869 7837 24903 7871
rect 20545 7769 20579 7803
rect 23857 7769 23891 7803
rect 18797 7701 18831 7735
rect 24685 7701 24719 7735
rect 21281 7429 21315 7463
rect 20269 7361 20303 7395
rect 22109 7361 22143 7395
rect 24133 7361 24167 7395
rect 22569 7293 22603 7327
rect 24777 7293 24811 7327
rect 24869 6817 24903 6851
rect 18245 6749 18279 6783
rect 19625 6749 19659 6783
rect 20821 6749 20855 6783
rect 22845 6749 22879 6783
rect 23857 6749 23891 6783
rect 18429 6681 18463 6715
rect 22017 6681 22051 6715
rect 24685 6681 24719 6715
rect 19441 6613 19475 6647
rect 19533 6409 19567 6443
rect 21281 6341 21315 6375
rect 19441 6273 19475 6307
rect 20085 6273 20119 6307
rect 22109 6273 22143 6307
rect 24133 6273 24167 6307
rect 22569 6205 22603 6239
rect 24777 6205 24811 6239
rect 19993 5865 20027 5899
rect 24777 5865 24811 5899
rect 21189 5729 21223 5763
rect 23029 5729 23063 5763
rect 20177 5661 20211 5695
rect 20729 5661 20763 5695
rect 22569 5661 22603 5695
rect 24685 5593 24719 5627
rect 16037 5185 16071 5219
rect 17877 5185 17911 5219
rect 19625 5185 19659 5219
rect 22017 5185 22051 5219
rect 24133 5185 24167 5219
rect 18981 5117 19015 5151
rect 20085 5117 20119 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 16129 4981 16163 5015
rect 25329 4777 25363 4811
rect 23489 4641 23523 4675
rect 17509 4573 17543 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 23213 4573 23247 4607
rect 18337 4505 18371 4539
rect 20361 4505 20395 4539
rect 22201 4505 22235 4539
rect 1777 4097 1811 4131
rect 7849 4097 7883 4131
rect 9321 4097 9355 4131
rect 13185 4097 13219 4131
rect 16865 4097 16899 4131
rect 18705 4097 18739 4131
rect 22109 4097 22143 4131
rect 23857 4097 23891 4131
rect 13461 4029 13495 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 24317 4029 24351 4063
rect 1593 3961 1627 3995
rect 8033 3961 8067 3995
rect 9505 3961 9539 3995
rect 2329 3689 2363 3723
rect 3249 3689 3283 3723
rect 5089 3689 5123 3723
rect 6561 3689 6595 3723
rect 7665 3689 7699 3723
rect 8401 3689 8435 3723
rect 9505 3689 9539 3723
rect 11529 3689 11563 3723
rect 1869 3621 1903 3655
rect 5641 3621 5675 3655
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 19901 3553 19935 3587
rect 23489 3553 23523 3587
rect 2513 3485 2547 3519
rect 3065 3485 3099 3519
rect 4905 3485 4939 3519
rect 5825 3485 5859 3519
rect 6377 3485 6411 3519
rect 7481 3485 7515 3519
rect 8217 3485 8251 3519
rect 9321 3485 9355 3519
rect 10057 3485 10091 3519
rect 10333 3485 10367 3519
rect 11345 3485 11379 3519
rect 12449 3485 12483 3519
rect 14289 3485 14323 3519
rect 16129 3485 16163 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 23213 3485 23247 3519
rect 1685 3417 1719 3451
rect 22201 3417 22235 3451
rect 2145 3145 2179 3179
rect 5181 3145 5215 3179
rect 24869 3145 24903 3179
rect 3065 3077 3099 3111
rect 6009 3077 6043 3111
rect 1961 3009 1995 3043
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 4261 3009 4295 3043
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 7389 3009 7423 3043
rect 8861 3009 8895 3043
rect 10609 3009 10643 3043
rect 11989 3009 12023 3043
rect 13001 3009 13035 3043
rect 14841 3009 14875 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 23581 3009 23615 3043
rect 7113 2941 7147 2975
rect 8585 2941 8619 2975
rect 10333 2941 10367 2975
rect 11713 2941 11747 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 22293 2941 22327 2975
rect 22569 2941 22603 2975
rect 3709 2873 3743 2907
rect 4445 2805 4479 2839
rect 2053 2601 2087 2635
rect 5917 2601 5951 2635
rect 11713 2601 11747 2635
rect 7297 2533 7331 2567
rect 4445 2465 4479 2499
rect 7757 2465 7791 2499
rect 14933 2465 14967 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 1869 2397 1903 2431
rect 2789 2397 2823 2431
rect 4169 2397 4203 2431
rect 5733 2397 5767 2431
rect 8033 2397 8067 2431
rect 9781 2397 9815 2431
rect 11897 2397 11931 2431
rect 12357 2397 12391 2431
rect 14657 2397 14691 2431
rect 16865 2397 16899 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 7113 2329 7147 2363
rect 10977 2329 11011 2363
rect 13277 2329 13311 2363
rect 2605 2261 2639 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 3237 54247 3295 54253
rect 3237 54213 3249 54247
rect 3283 54244 3295 54247
rect 5350 54244 5356 54256
rect 3283 54216 5356 54244
rect 3283 54213 3295 54216
rect 3237 54207 3295 54213
rect 5350 54204 5356 54216
rect 5408 54204 5414 54256
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 6822 54244 6828 54256
rect 5859 54216 6828 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 6822 54204 6828 54216
rect 6880 54204 6886 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 9398 54244 9404 54256
rect 8435 54216 9404 54244
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 9398 54204 9404 54216
rect 9456 54204 9462 54256
rect 10870 54204 10876 54256
rect 10928 54204 10934 54256
rect 14918 54204 14924 54256
rect 14976 54244 14982 54256
rect 15473 54247 15531 54253
rect 15473 54244 15485 54247
rect 14976 54216 15485 54244
rect 14976 54204 14982 54216
rect 15473 54213 15485 54216
rect 15519 54213 15531 54247
rect 15473 54207 15531 54213
rect 16022 54204 16028 54256
rect 16080 54244 16086 54256
rect 16080 54216 16574 54244
rect 16080 54204 16086 54216
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4706 54176 4712 54188
rect 2271 54148 4712 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4706 54136 4712 54148
rect 4764 54136 4770 54188
rect 4801 54179 4859 54185
rect 4801 54145 4813 54179
rect 4847 54176 4859 54179
rect 7377 54179 7435 54185
rect 4847 54148 6914 54176
rect 4847 54145 4859 54148
rect 4801 54139 4859 54145
rect 6886 54108 6914 54148
rect 7377 54145 7389 54179
rect 7423 54176 7435 54179
rect 7466 54176 7472 54188
rect 7423 54148 7472 54176
rect 7423 54145 7435 54148
rect 7377 54139 7435 54145
rect 7466 54136 7472 54148
rect 7524 54136 7530 54188
rect 9858 54136 9864 54188
rect 9916 54136 9922 54188
rect 12066 54136 12072 54188
rect 12124 54136 12130 54188
rect 14550 54136 14556 54188
rect 14608 54176 14614 54188
rect 14645 54179 14703 54185
rect 14645 54176 14657 54179
rect 14608 54148 14657 54176
rect 14608 54136 14614 54148
rect 14645 54145 14657 54148
rect 14691 54145 14703 54179
rect 14645 54139 14703 54145
rect 15286 54136 15292 54188
rect 15344 54176 15350 54188
rect 16301 54179 16359 54185
rect 16301 54176 16313 54179
rect 15344 54148 16313 54176
rect 15344 54136 15350 54148
rect 16301 54145 16313 54148
rect 16347 54145 16359 54179
rect 16546 54176 16574 54216
rect 17126 54204 17132 54256
rect 17184 54244 17190 54256
rect 17681 54247 17739 54253
rect 17681 54244 17693 54247
rect 17184 54216 17693 54244
rect 17184 54204 17190 54216
rect 17681 54213 17693 54216
rect 17727 54213 17739 54247
rect 17681 54207 17739 54213
rect 19334 54204 19340 54256
rect 19392 54244 19398 54256
rect 19392 54216 19564 54244
rect 19392 54204 19398 54216
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 16301 54139 16359 54145
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 17494 54136 17500 54188
rect 17552 54176 17558 54188
rect 18417 54179 18475 54185
rect 18417 54176 18429 54179
rect 17552 54148 18429 54176
rect 17552 54136 17558 54148
rect 18417 54145 18429 54148
rect 18463 54145 18475 54179
rect 18417 54139 18475 54145
rect 18598 54136 18604 54188
rect 18656 54176 18662 54188
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 18656 54148 19441 54176
rect 18656 54136 18662 54148
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19536 54176 19564 54216
rect 20070 54204 20076 54256
rect 20128 54244 20134 54256
rect 23845 54247 23903 54253
rect 20128 54216 20944 54244
rect 20128 54204 20134 54216
rect 20916 54185 20944 54216
rect 23845 54213 23857 54247
rect 23891 54244 23903 54247
rect 24118 54244 24124 54256
rect 23891 54216 24124 54244
rect 23891 54213 23903 54216
rect 23845 54207 23903 54213
rect 24118 54204 24124 54216
rect 24176 54204 24182 54256
rect 20257 54179 20315 54185
rect 20257 54176 20269 54179
rect 19536 54148 20269 54176
rect 19429 54139 19487 54145
rect 20257 54145 20269 54148
rect 20303 54145 20315 54179
rect 20257 54139 20315 54145
rect 20901 54179 20959 54185
rect 20901 54145 20913 54179
rect 20947 54145 20959 54179
rect 20901 54139 20959 54145
rect 21174 54136 21180 54188
rect 21232 54176 21238 54188
rect 22189 54179 22247 54185
rect 22189 54176 22201 54179
rect 21232 54148 22201 54176
rect 21232 54136 21238 54148
rect 22189 54145 22201 54148
rect 22235 54145 22247 54179
rect 22189 54139 22247 54145
rect 22649 54179 22707 54185
rect 22649 54145 22661 54179
rect 22695 54145 22707 54179
rect 22649 54139 22707 54145
rect 8570 54108 8576 54120
rect 6886 54080 8576 54108
rect 8570 54068 8576 54080
rect 8628 54068 8634 54120
rect 11974 54068 11980 54120
rect 12032 54108 12038 54120
rect 12529 54111 12587 54117
rect 12529 54108 12541 54111
rect 12032 54080 12541 54108
rect 12032 54068 12038 54080
rect 12529 54077 12541 54080
rect 12575 54077 12587 54111
rect 22664 54108 22692 54139
rect 22738 54136 22744 54188
rect 22796 54176 22802 54188
rect 24765 54179 24823 54185
rect 24765 54176 24777 54179
rect 22796 54148 24777 54176
rect 22796 54136 22802 54148
rect 24765 54145 24777 54148
rect 24811 54145 24823 54179
rect 24765 54139 24823 54145
rect 23750 54108 23756 54120
rect 22664 54080 23756 54108
rect 12529 54071 12587 54077
rect 23750 54068 23756 54080
rect 23808 54068 23814 54120
rect 15746 54000 15752 54052
rect 15804 54040 15810 54052
rect 17037 54043 17095 54049
rect 17037 54040 17049 54043
rect 15804 54012 17049 54040
rect 15804 54000 15810 54012
rect 17037 54009 17049 54012
rect 17083 54009 17095 54043
rect 17037 54003 17095 54009
rect 20441 54043 20499 54049
rect 20441 54009 20453 54043
rect 20487 54040 20499 54043
rect 20622 54040 20628 54052
rect 20487 54012 20628 54040
rect 20487 54009 20499 54012
rect 20441 54003 20499 54009
rect 20622 54000 20628 54012
rect 20680 54000 20686 54052
rect 14826 53932 14832 53984
rect 14884 53932 14890 53984
rect 15562 53932 15568 53984
rect 15620 53932 15626 53984
rect 16114 53932 16120 53984
rect 16172 53932 16178 53984
rect 17770 53932 17776 53984
rect 17828 53932 17834 53984
rect 18506 53932 18512 53984
rect 18564 53932 18570 53984
rect 19610 53932 19616 53984
rect 19668 53932 19674 53984
rect 20990 53932 20996 53984
rect 21048 53972 21054 53984
rect 21085 53975 21143 53981
rect 21085 53972 21097 53975
rect 21048 53944 21097 53972
rect 21048 53932 21054 53944
rect 21085 53941 21097 53944
rect 21131 53941 21143 53975
rect 21085 53935 21143 53941
rect 21818 53932 21824 53984
rect 21876 53972 21882 53984
rect 22005 53975 22063 53981
rect 22005 53972 22017 53975
rect 21876 53944 22017 53972
rect 21876 53932 21882 53944
rect 22005 53941 22017 53944
rect 22051 53941 22063 53975
rect 22005 53935 22063 53941
rect 23382 53932 23388 53984
rect 23440 53972 23446 53984
rect 24581 53975 24639 53981
rect 24581 53972 24593 53975
rect 23440 53944 24593 53972
rect 23440 53932 23446 53944
rect 24581 53941 24593 53944
rect 24627 53941 24639 53975
rect 24581 53935 24639 53941
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 3237 53635 3295 53641
rect 3237 53601 3249 53635
rect 3283 53632 3295 53635
rect 4614 53632 4620 53644
rect 3283 53604 4620 53632
rect 3283 53601 3295 53604
rect 3237 53595 3295 53601
rect 4614 53592 4620 53604
rect 4672 53592 4678 53644
rect 6549 53635 6607 53641
rect 6549 53601 6561 53635
rect 6595 53632 6607 53635
rect 7558 53632 7564 53644
rect 6595 53604 7564 53632
rect 6595 53601 6607 53604
rect 6549 53595 6607 53601
rect 7558 53592 7564 53604
rect 7616 53592 7622 53644
rect 8294 53592 8300 53644
rect 8352 53592 8358 53644
rect 9030 53592 9036 53644
rect 9088 53632 9094 53644
rect 9674 53632 9680 53644
rect 9088 53604 9680 53632
rect 9088 53592 9094 53604
rect 9674 53592 9680 53604
rect 9732 53592 9738 53644
rect 10502 53592 10508 53644
rect 10560 53592 10566 53644
rect 11606 53592 11612 53644
rect 11664 53632 11670 53644
rect 12161 53635 12219 53641
rect 12161 53632 12173 53635
rect 11664 53604 12173 53632
rect 11664 53592 11670 53604
rect 12161 53601 12173 53604
rect 12207 53601 12219 53635
rect 12161 53595 12219 53601
rect 23845 53635 23903 53641
rect 23845 53601 23857 53635
rect 23891 53632 23903 53635
rect 25590 53632 25596 53644
rect 23891 53604 25596 53632
rect 23891 53601 23903 53604
rect 23845 53595 23903 53601
rect 25590 53592 25596 53604
rect 25648 53592 25654 53644
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53533 2283 53567
rect 2225 53527 2283 53533
rect 2240 53496 2268 53527
rect 5442 53524 5448 53576
rect 5500 53524 5506 53576
rect 7374 53524 7380 53576
rect 7432 53524 7438 53576
rect 10042 53524 10048 53576
rect 10100 53524 10106 53576
rect 11698 53524 11704 53576
rect 11756 53524 11762 53576
rect 13725 53567 13783 53573
rect 13725 53533 13737 53567
rect 13771 53564 13783 53567
rect 13814 53564 13820 53576
rect 13771 53536 13820 53564
rect 13771 53533 13783 53536
rect 13725 53527 13783 53533
rect 13814 53524 13820 53536
rect 13872 53524 13878 53576
rect 14182 53524 14188 53576
rect 14240 53564 14246 53576
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 14240 53536 14289 53564
rect 14240 53524 14246 53536
rect 14277 53533 14289 53536
rect 14323 53533 14335 53567
rect 14277 53527 14335 53533
rect 15654 53524 15660 53576
rect 15712 53564 15718 53576
rect 15749 53567 15807 53573
rect 15749 53564 15761 53567
rect 15712 53536 15761 53564
rect 15712 53524 15718 53536
rect 15749 53533 15761 53536
rect 15795 53533 15807 53567
rect 15749 53527 15807 53533
rect 16390 53524 16396 53576
rect 16448 53564 16454 53576
rect 16485 53567 16543 53573
rect 16485 53564 16497 53567
rect 16448 53536 16497 53564
rect 16448 53524 16454 53536
rect 16485 53533 16497 53536
rect 16531 53533 16543 53567
rect 16485 53527 16543 53533
rect 16758 53524 16764 53576
rect 16816 53564 16822 53576
rect 17405 53567 17463 53573
rect 17405 53564 17417 53567
rect 16816 53536 17417 53564
rect 16816 53524 16822 53536
rect 17405 53533 17417 53536
rect 17451 53533 17463 53567
rect 17405 53527 17463 53533
rect 17862 53524 17868 53576
rect 17920 53564 17926 53576
rect 18049 53567 18107 53573
rect 18049 53564 18061 53567
rect 17920 53536 18061 53564
rect 17920 53524 17926 53536
rect 18049 53533 18061 53536
rect 18095 53533 18107 53567
rect 18049 53527 18107 53533
rect 18322 53524 18328 53576
rect 18380 53564 18386 53576
rect 18877 53567 18935 53573
rect 18877 53564 18889 53567
rect 18380 53536 18889 53564
rect 18380 53524 18386 53536
rect 18877 53533 18889 53536
rect 18923 53533 18935 53567
rect 18877 53527 18935 53533
rect 18966 53524 18972 53576
rect 19024 53564 19030 53576
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 19024 53536 19441 53564
rect 19024 53524 19030 53536
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 20438 53524 20444 53576
rect 20496 53564 20502 53576
rect 20533 53567 20591 53573
rect 20533 53564 20545 53567
rect 20496 53536 20545 53564
rect 20496 53524 20502 53536
rect 20533 53533 20545 53536
rect 20579 53533 20591 53567
rect 20533 53527 20591 53533
rect 20806 53524 20812 53576
rect 20864 53564 20870 53576
rect 21269 53567 21327 53573
rect 21269 53564 21281 53567
rect 20864 53536 21281 53564
rect 20864 53524 20870 53536
rect 21269 53533 21281 53536
rect 21315 53533 21327 53567
rect 21269 53527 21327 53533
rect 21542 53524 21548 53576
rect 21600 53564 21606 53576
rect 22189 53567 22247 53573
rect 22189 53564 22201 53567
rect 21600 53536 22201 53564
rect 21600 53524 21606 53536
rect 22189 53533 22201 53536
rect 22235 53533 22247 53567
rect 22189 53527 22247 53533
rect 22833 53567 22891 53573
rect 22833 53533 22845 53567
rect 22879 53533 22891 53567
rect 22833 53527 22891 53533
rect 6638 53496 6644 53508
rect 2240 53468 6644 53496
rect 6638 53456 6644 53468
rect 6696 53456 6702 53508
rect 18233 53499 18291 53505
rect 18233 53465 18245 53499
rect 18279 53496 18291 53499
rect 18414 53496 18420 53508
rect 18279 53468 18420 53496
rect 18279 53465 18291 53468
rect 18233 53459 18291 53465
rect 18414 53456 18420 53468
rect 18472 53456 18478 53508
rect 22848 53496 22876 53527
rect 23290 53524 23296 53576
rect 23348 53564 23354 53576
rect 24765 53567 24823 53573
rect 24765 53564 24777 53567
rect 23348 53536 24777 53564
rect 23348 53524 23354 53536
rect 24765 53533 24777 53536
rect 24811 53533 24823 53567
rect 24765 53527 24823 53533
rect 25866 53496 25872 53508
rect 20732 53468 21588 53496
rect 22848 53468 25872 53496
rect 12526 53388 12532 53440
rect 12584 53428 12590 53440
rect 13541 53431 13599 53437
rect 13541 53428 13553 53431
rect 12584 53400 13553 53428
rect 12584 53388 12590 53400
rect 13541 53397 13553 53400
rect 13587 53397 13599 53431
rect 13541 53391 13599 53397
rect 14458 53388 14464 53440
rect 14516 53388 14522 53440
rect 15930 53388 15936 53440
rect 15988 53388 15994 53440
rect 16206 53388 16212 53440
rect 16264 53428 16270 53440
rect 16669 53431 16727 53437
rect 16669 53428 16681 53431
rect 16264 53400 16681 53428
rect 16264 53388 16270 53400
rect 16669 53397 16681 53400
rect 16715 53397 16727 53431
rect 16669 53391 16727 53397
rect 17218 53388 17224 53440
rect 17276 53388 17282 53440
rect 18690 53388 18696 53440
rect 18748 53388 18754 53440
rect 19613 53431 19671 53437
rect 19613 53397 19625 53431
rect 19659 53428 19671 53431
rect 20070 53428 20076 53440
rect 19659 53400 20076 53428
rect 19659 53397 19671 53400
rect 19613 53391 19671 53397
rect 20070 53388 20076 53400
rect 20128 53388 20134 53440
rect 20732 53437 20760 53468
rect 21560 53440 21588 53468
rect 25866 53456 25872 53468
rect 25924 53456 25930 53508
rect 20717 53431 20775 53437
rect 20717 53397 20729 53431
rect 20763 53397 20775 53431
rect 20717 53391 20775 53397
rect 21450 53388 21456 53440
rect 21508 53388 21514 53440
rect 21542 53388 21548 53440
rect 21600 53388 21606 53440
rect 22002 53388 22008 53440
rect 22060 53388 22066 53440
rect 23290 53388 23296 53440
rect 23348 53428 23354 53440
rect 24581 53431 24639 53437
rect 24581 53428 24593 53431
rect 23348 53400 24593 53428
rect 23348 53388 23354 53400
rect 24581 53397 24593 53400
rect 24627 53397 24639 53431
rect 24581 53391 24639 53397
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 2774 53224 2780 53236
rect 1780 53196 2780 53224
rect 1780 53097 1808 53196
rect 2774 53184 2780 53196
rect 2832 53184 2838 53236
rect 3973 53159 4031 53165
rect 3973 53125 3985 53159
rect 4019 53156 4031 53159
rect 4246 53156 4252 53168
rect 4019 53128 4252 53156
rect 4019 53125 4031 53128
rect 3973 53119 4031 53125
rect 4246 53116 4252 53128
rect 4304 53116 4310 53168
rect 5718 53116 5724 53168
rect 5776 53116 5782 53168
rect 12710 53116 12716 53168
rect 12768 53156 12774 53168
rect 14369 53159 14427 53165
rect 14369 53156 14381 53159
rect 12768 53128 14381 53156
rect 12768 53116 12774 53128
rect 14369 53125 14381 53128
rect 14415 53125 14427 53159
rect 14369 53119 14427 53125
rect 24854 53116 24860 53168
rect 24912 53116 24918 53168
rect 1765 53091 1823 53097
rect 1765 53057 1777 53091
rect 1811 53057 1823 53091
rect 1765 53051 1823 53057
rect 2961 53091 3019 53097
rect 2961 53057 2973 53091
rect 3007 53057 3019 53091
rect 2961 53051 3019 53057
rect 4801 53091 4859 53097
rect 4801 53057 4813 53091
rect 4847 53088 4859 53091
rect 6362 53088 6368 53100
rect 4847 53060 6368 53088
rect 4847 53057 4859 53060
rect 4801 53051 4859 53057
rect 2976 53020 3004 53051
rect 6362 53048 6368 53060
rect 6420 53048 6426 53100
rect 6822 53048 6828 53100
rect 6880 53048 6886 53100
rect 8113 53091 8171 53097
rect 8113 53057 8125 53091
rect 8159 53088 8171 53091
rect 9214 53088 9220 53100
rect 8159 53060 9220 53088
rect 8159 53057 8171 53060
rect 8113 53051 8171 53057
rect 9214 53048 9220 53060
rect 9272 53048 9278 53100
rect 9398 53048 9404 53100
rect 9456 53088 9462 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9456 53060 9781 53088
rect 9456 53048 9462 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 10502 53048 10508 53100
rect 10560 53088 10566 53100
rect 11701 53091 11759 53097
rect 11701 53088 11713 53091
rect 10560 53060 11713 53088
rect 10560 53048 10566 53060
rect 11701 53057 11713 53060
rect 11747 53057 11759 53091
rect 11701 53051 11759 53057
rect 13446 53048 13452 53100
rect 13504 53088 13510 53100
rect 13541 53091 13599 53097
rect 13541 53088 13553 53091
rect 13504 53060 13553 53088
rect 13504 53048 13510 53060
rect 13541 53057 13553 53060
rect 13587 53057 13599 53091
rect 13541 53051 13599 53057
rect 19702 53048 19708 53100
rect 19760 53088 19766 53100
rect 19981 53091 20039 53097
rect 19981 53088 19993 53091
rect 19760 53060 19993 53088
rect 19760 53048 19766 53060
rect 19981 53057 19993 53060
rect 20027 53057 20039 53091
rect 19981 53051 20039 53057
rect 21910 53048 21916 53100
rect 21968 53088 21974 53100
rect 22005 53091 22063 53097
rect 22005 53088 22017 53091
rect 21968 53060 22017 53088
rect 21968 53048 21974 53060
rect 22005 53057 22017 53060
rect 22051 53057 22063 53091
rect 22005 53051 22063 53057
rect 22278 53048 22284 53100
rect 22336 53088 22342 53100
rect 22925 53091 22983 53097
rect 22925 53088 22937 53091
rect 22336 53060 22937 53088
rect 22336 53048 22342 53060
rect 22925 53057 22937 53060
rect 22971 53057 22983 53091
rect 22925 53051 22983 53057
rect 24121 53091 24179 53097
rect 24121 53057 24133 53091
rect 24167 53088 24179 53091
rect 25958 53088 25964 53100
rect 24167 53060 25964 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 25958 53048 25964 53060
rect 26016 53048 26022 53100
rect 6546 53020 6552 53032
rect 2976 52992 6552 53020
rect 6546 52980 6552 52992
rect 6604 52980 6610 53032
rect 8662 52980 8668 53032
rect 8720 52980 8726 53032
rect 10134 52980 10140 53032
rect 10192 53020 10198 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10192 52992 10241 53020
rect 10192 52980 10198 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 11238 52980 11244 53032
rect 11296 53020 11302 53032
rect 12161 53023 12219 53029
rect 12161 53020 12173 53023
rect 11296 52992 12173 53020
rect 11296 52980 11302 52992
rect 12161 52989 12173 52992
rect 12207 52989 12219 53023
rect 12161 52983 12219 52989
rect 14550 52912 14556 52964
rect 14608 52912 14614 52964
rect 1581 52887 1639 52893
rect 1581 52853 1593 52887
rect 1627 52884 1639 52887
rect 3970 52884 3976 52896
rect 1627 52856 3976 52884
rect 1627 52853 1639 52856
rect 1581 52847 1639 52853
rect 3970 52844 3976 52856
rect 4028 52844 4034 52896
rect 4246 52844 4252 52896
rect 4304 52884 4310 52896
rect 6641 52887 6699 52893
rect 6641 52884 6653 52887
rect 4304 52856 6653 52884
rect 4304 52844 4310 52856
rect 6641 52853 6653 52856
rect 6687 52853 6699 52887
rect 6641 52847 6699 52853
rect 13722 52844 13728 52896
rect 13780 52844 13786 52896
rect 19794 52844 19800 52896
rect 19852 52844 19858 52896
rect 22186 52844 22192 52896
rect 22244 52844 22250 52896
rect 22738 52844 22744 52896
rect 22796 52844 22802 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 2038 52640 2044 52692
rect 2096 52680 2102 52692
rect 3418 52680 3424 52692
rect 2096 52652 3424 52680
rect 2096 52640 2102 52652
rect 3418 52640 3424 52652
rect 3476 52640 3482 52692
rect 11793 52683 11851 52689
rect 11793 52649 11805 52683
rect 11839 52680 11851 52683
rect 12066 52680 12072 52692
rect 11839 52652 12072 52680
rect 11839 52649 11851 52652
rect 11793 52643 11851 52649
rect 12066 52640 12072 52652
rect 12124 52640 12130 52692
rect 23750 52640 23756 52692
rect 23808 52640 23814 52692
rect 934 52572 940 52624
rect 992 52612 998 52624
rect 4430 52612 4436 52624
rect 992 52584 4436 52612
rect 992 52572 998 52584
rect 4430 52572 4436 52584
rect 4488 52572 4494 52624
rect 12437 52615 12495 52621
rect 12437 52581 12449 52615
rect 12483 52612 12495 52615
rect 13446 52612 13452 52624
rect 12483 52584 13452 52612
rect 12483 52581 12495 52584
rect 12437 52575 12495 52581
rect 13446 52572 13452 52584
rect 13504 52572 13510 52624
rect 1302 52504 1308 52556
rect 1360 52544 1366 52556
rect 3973 52547 4031 52553
rect 3973 52544 3985 52547
rect 1360 52516 3985 52544
rect 1360 52504 1366 52516
rect 3973 52513 3985 52516
rect 4019 52513 4031 52547
rect 3973 52507 4031 52513
rect 4249 52547 4307 52553
rect 4249 52513 4261 52547
rect 4295 52544 4307 52547
rect 5994 52544 6000 52556
rect 4295 52516 6000 52544
rect 4295 52513 4307 52516
rect 4249 52507 4307 52513
rect 5994 52504 6000 52516
rect 6052 52504 6058 52556
rect 6086 52504 6092 52556
rect 6144 52504 6150 52556
rect 7834 52504 7840 52556
rect 7892 52504 7898 52556
rect 9766 52504 9772 52556
rect 9824 52544 9830 52556
rect 10321 52547 10379 52553
rect 10321 52544 10333 52547
rect 9824 52516 10333 52544
rect 9824 52504 9830 52516
rect 10321 52513 10333 52516
rect 10367 52513 10379 52547
rect 10321 52507 10379 52513
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 3142 52476 3148 52488
rect 2271 52448 3148 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 3142 52436 3148 52448
rect 3200 52436 3206 52488
rect 3237 52479 3295 52485
rect 3237 52445 3249 52479
rect 3283 52476 3295 52479
rect 3326 52476 3332 52488
rect 3283 52448 3332 52476
rect 3283 52445 3295 52448
rect 3237 52439 3295 52445
rect 3326 52436 3332 52448
rect 3384 52436 3390 52488
rect 5445 52479 5503 52485
rect 5445 52445 5457 52479
rect 5491 52476 5503 52479
rect 5718 52476 5724 52488
rect 5491 52448 5724 52476
rect 5491 52445 5503 52448
rect 5445 52439 5503 52445
rect 5718 52436 5724 52448
rect 5776 52436 5782 52488
rect 6454 52436 6460 52488
rect 6512 52476 6518 52488
rect 6914 52476 6920 52488
rect 6512 52448 6920 52476
rect 6512 52436 6518 52448
rect 6914 52436 6920 52448
rect 6972 52436 6978 52488
rect 7377 52479 7435 52485
rect 7377 52445 7389 52479
rect 7423 52476 7435 52479
rect 8938 52476 8944 52488
rect 7423 52448 8944 52476
rect 7423 52445 7435 52448
rect 7377 52439 7435 52445
rect 8938 52436 8944 52448
rect 8996 52436 9002 52488
rect 9582 52436 9588 52488
rect 9640 52476 9646 52488
rect 9861 52479 9919 52485
rect 9861 52476 9873 52479
rect 9640 52448 9873 52476
rect 9640 52436 9646 52448
rect 9861 52445 9873 52448
rect 9907 52445 9919 52479
rect 9861 52439 9919 52445
rect 11974 52436 11980 52488
rect 12032 52436 12038 52488
rect 12342 52436 12348 52488
rect 12400 52476 12406 52488
rect 12621 52479 12679 52485
rect 12621 52476 12633 52479
rect 12400 52448 12633 52476
rect 12400 52436 12406 52448
rect 12621 52445 12633 52448
rect 12667 52445 12679 52479
rect 12621 52439 12679 52445
rect 13354 52436 13360 52488
rect 13412 52436 13418 52488
rect 13449 52479 13507 52485
rect 13449 52445 13461 52479
rect 13495 52476 13507 52479
rect 14090 52476 14096 52488
rect 13495 52448 14096 52476
rect 13495 52445 13507 52448
rect 13449 52439 13507 52445
rect 14090 52436 14096 52448
rect 14148 52436 14154 52488
rect 23937 52479 23995 52485
rect 23937 52445 23949 52479
rect 23983 52476 23995 52479
rect 24486 52476 24492 52488
rect 23983 52448 24492 52476
rect 23983 52445 23995 52448
rect 23937 52439 23995 52445
rect 24486 52436 24492 52448
rect 24544 52436 24550 52488
rect 13265 52411 13323 52417
rect 13265 52377 13277 52411
rect 13311 52408 13323 52411
rect 13372 52408 13400 52436
rect 13311 52380 13400 52408
rect 13311 52377 13323 52380
rect 13265 52371 13323 52377
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 11698 52096 11704 52148
rect 11756 52096 11762 52148
rect 5626 52068 5632 52080
rect 2976 52040 5632 52068
rect 2976 52009 3004 52040
rect 5626 52028 5632 52040
rect 5684 52028 5690 52080
rect 2961 52003 3019 52009
rect 2961 51969 2973 52003
rect 3007 51969 3019 52003
rect 2961 51963 3019 51969
rect 4801 52003 4859 52009
rect 4801 51969 4813 52003
rect 4847 52000 4859 52003
rect 6270 52000 6276 52012
rect 4847 51972 6276 52000
rect 4847 51969 4859 51972
rect 4801 51963 4859 51969
rect 6270 51960 6276 51972
rect 6328 51960 6334 52012
rect 7098 51960 7104 52012
rect 7156 51960 7162 52012
rect 9122 51960 9128 52012
rect 9180 51960 9186 52012
rect 11882 51960 11888 52012
rect 11940 51960 11946 52012
rect 25130 51960 25136 52012
rect 25188 51960 25194 52012
rect 3510 51892 3516 51944
rect 3568 51892 3574 51944
rect 4982 51892 4988 51944
rect 5040 51932 5046 51944
rect 5077 51935 5135 51941
rect 5077 51932 5089 51935
rect 5040 51904 5089 51932
rect 5040 51892 5046 51904
rect 5077 51901 5089 51904
rect 5123 51901 5135 51935
rect 5077 51895 5135 51901
rect 7006 51892 7012 51944
rect 7064 51932 7070 51944
rect 7377 51935 7435 51941
rect 7377 51932 7389 51935
rect 7064 51904 7389 51932
rect 7064 51892 7070 51904
rect 7377 51901 7389 51904
rect 7423 51901 7435 51935
rect 7377 51895 7435 51901
rect 9674 51892 9680 51944
rect 9732 51892 9738 51944
rect 24118 51756 24124 51808
rect 24176 51796 24182 51808
rect 25225 51799 25283 51805
rect 25225 51796 25237 51799
rect 24176 51768 25237 51796
rect 24176 51756 24182 51768
rect 25225 51765 25237 51768
rect 25271 51765 25283 51799
rect 25225 51759 25283 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 4706 51552 4712 51604
rect 4764 51592 4770 51604
rect 5905 51595 5963 51601
rect 5905 51592 5917 51595
rect 4764 51564 5917 51592
rect 4764 51552 4770 51564
rect 5905 51561 5917 51564
rect 5951 51561 5963 51595
rect 5905 51555 5963 51561
rect 2774 51416 2780 51468
rect 2832 51416 2838 51468
rect 4154 51416 4160 51468
rect 4212 51456 4218 51468
rect 4433 51459 4491 51465
rect 4433 51456 4445 51459
rect 4212 51428 4445 51456
rect 4212 51416 4218 51428
rect 4433 51425 4445 51428
rect 4479 51425 4491 51459
rect 4433 51419 4491 51425
rect 6914 51416 6920 51468
rect 6972 51456 6978 51468
rect 7009 51459 7067 51465
rect 7009 51456 7021 51459
rect 6972 51428 7021 51456
rect 6972 51416 6978 51428
rect 7009 51425 7021 51428
rect 7055 51425 7067 51459
rect 7009 51419 7067 51425
rect 2225 51391 2283 51397
rect 2225 51357 2237 51391
rect 2271 51357 2283 51391
rect 2225 51351 2283 51357
rect 4065 51391 4123 51397
rect 4065 51357 4077 51391
rect 4111 51388 4123 51391
rect 4246 51388 4252 51400
rect 4111 51360 4252 51388
rect 4111 51357 4123 51360
rect 4065 51351 4123 51357
rect 2240 51252 2268 51351
rect 4246 51348 4252 51360
rect 4304 51348 4310 51400
rect 6089 51391 6147 51397
rect 6089 51357 6101 51391
rect 6135 51357 6147 51391
rect 6089 51351 6147 51357
rect 6733 51391 6791 51397
rect 6733 51357 6745 51391
rect 6779 51388 6791 51391
rect 7282 51388 7288 51400
rect 6779 51360 7288 51388
rect 6779 51357 6791 51360
rect 6733 51351 6791 51357
rect 6104 51320 6132 51351
rect 7282 51348 7288 51360
rect 7340 51348 7346 51400
rect 25038 51348 25044 51400
rect 25096 51348 25102 51400
rect 7006 51320 7012 51332
rect 6104 51292 7012 51320
rect 7006 51280 7012 51292
rect 7064 51280 7070 51332
rect 5534 51252 5540 51264
rect 2240 51224 5540 51252
rect 5534 51212 5540 51224
rect 5592 51212 5598 51264
rect 25225 51255 25283 51261
rect 25225 51221 25237 51255
rect 25271 51252 25283 51255
rect 25590 51252 25596 51264
rect 25271 51224 25596 51252
rect 25271 51221 25283 51224
rect 25225 51215 25283 51221
rect 25590 51212 25596 51224
rect 25648 51212 25654 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 5534 51008 5540 51060
rect 5592 51048 5598 51060
rect 6917 51051 6975 51057
rect 6917 51048 6929 51051
rect 5592 51020 6929 51048
rect 5592 51008 5598 51020
rect 6917 51017 6929 51020
rect 6963 51017 6975 51051
rect 6917 51011 6975 51017
rect 9858 51008 9864 51060
rect 9916 51008 9922 51060
rect 10502 51008 10508 51060
rect 10560 51008 10566 51060
rect 3053 50915 3111 50921
rect 3053 50881 3065 50915
rect 3099 50912 3111 50915
rect 3694 50912 3700 50924
rect 3099 50884 3700 50912
rect 3099 50881 3111 50884
rect 3053 50875 3111 50881
rect 3694 50872 3700 50884
rect 3752 50872 3758 50924
rect 6825 50915 6883 50921
rect 6825 50881 6837 50915
rect 6871 50912 6883 50915
rect 7190 50912 7196 50924
rect 6871 50884 7196 50912
rect 6871 50881 6883 50884
rect 6825 50875 6883 50881
rect 7190 50872 7196 50884
rect 7248 50872 7254 50924
rect 8386 50872 8392 50924
rect 8444 50912 8450 50924
rect 9769 50915 9827 50921
rect 9769 50912 9781 50915
rect 8444 50884 9781 50912
rect 8444 50872 8450 50884
rect 9769 50881 9781 50884
rect 9815 50881 9827 50915
rect 9769 50875 9827 50881
rect 9950 50872 9956 50924
rect 10008 50912 10014 50924
rect 10689 50915 10747 50921
rect 10689 50912 10701 50915
rect 10008 50884 10701 50912
rect 10008 50872 10014 50884
rect 10689 50881 10701 50884
rect 10735 50881 10747 50915
rect 10689 50875 10747 50881
rect 25038 50872 25044 50924
rect 25096 50872 25102 50924
rect 934 50804 940 50856
rect 992 50844 998 50856
rect 1581 50847 1639 50853
rect 1581 50844 1593 50847
rect 992 50816 1593 50844
rect 992 50804 998 50816
rect 1581 50813 1593 50816
rect 1627 50813 1639 50847
rect 1581 50807 1639 50813
rect 1857 50847 1915 50853
rect 1857 50813 1869 50847
rect 1903 50813 1915 50847
rect 1857 50807 1915 50813
rect 1872 50776 1900 50807
rect 2866 50804 2872 50856
rect 2924 50844 2930 50856
rect 3329 50847 3387 50853
rect 3329 50844 3341 50847
rect 2924 50816 3341 50844
rect 2924 50804 2930 50816
rect 3329 50813 3341 50816
rect 3375 50813 3387 50847
rect 3329 50807 3387 50813
rect 7558 50776 7564 50788
rect 1872 50748 7564 50776
rect 7558 50736 7564 50748
rect 7616 50736 7622 50788
rect 25225 50711 25283 50717
rect 25225 50677 25237 50711
rect 25271 50708 25283 50711
rect 25682 50708 25688 50720
rect 25271 50680 25688 50708
rect 25271 50677 25283 50680
rect 25225 50671 25283 50677
rect 25682 50668 25688 50680
rect 25740 50668 25746 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 6181 50507 6239 50513
rect 6181 50473 6193 50507
rect 6227 50504 6239 50507
rect 7098 50504 7104 50516
rect 6227 50476 7104 50504
rect 6227 50473 6239 50476
rect 6181 50467 6239 50473
rect 7098 50464 7104 50476
rect 7156 50464 7162 50516
rect 9398 50396 9404 50448
rect 9456 50396 9462 50448
rect 3237 50371 3295 50377
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 3418 50368 3424 50380
rect 3283 50340 3424 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 3418 50328 3424 50340
rect 3476 50328 3482 50380
rect 4430 50328 4436 50380
rect 4488 50328 4494 50380
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50300 2283 50303
rect 3510 50300 3516 50312
rect 2271 50272 3516 50300
rect 2271 50269 2283 50272
rect 2225 50263 2283 50269
rect 3510 50260 3516 50272
rect 3568 50260 3574 50312
rect 4065 50303 4123 50309
rect 4065 50269 4077 50303
rect 4111 50300 4123 50303
rect 4111 50272 5488 50300
rect 4111 50269 4123 50272
rect 4065 50263 4123 50269
rect 5460 50232 5488 50272
rect 5534 50260 5540 50312
rect 5592 50300 5598 50312
rect 6365 50303 6423 50309
rect 6365 50300 6377 50303
rect 5592 50272 6377 50300
rect 5592 50260 5598 50272
rect 6365 50269 6377 50272
rect 6411 50269 6423 50303
rect 6365 50263 6423 50269
rect 6914 50260 6920 50312
rect 6972 50300 6978 50312
rect 9217 50303 9275 50309
rect 9217 50300 9229 50303
rect 6972 50272 9229 50300
rect 6972 50260 6978 50272
rect 9217 50269 9229 50272
rect 9263 50269 9275 50303
rect 9217 50263 9275 50269
rect 25038 50260 25044 50312
rect 25096 50260 25102 50312
rect 10410 50232 10416 50244
rect 5460 50204 10416 50232
rect 10410 50192 10416 50204
rect 10468 50192 10474 50244
rect 25225 50167 25283 50173
rect 25225 50133 25237 50167
rect 25271 50164 25283 50167
rect 25774 50164 25780 50176
rect 25271 50136 25780 50164
rect 25271 50133 25283 50136
rect 25225 50127 25283 50133
rect 25774 50124 25780 50136
rect 25832 50124 25838 50176
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 7374 49920 7380 49972
rect 7432 49960 7438 49972
rect 7837 49963 7895 49969
rect 7837 49960 7849 49963
rect 7432 49932 7849 49960
rect 7432 49920 7438 49932
rect 7837 49929 7849 49932
rect 7883 49929 7895 49963
rect 7837 49923 7895 49929
rect 9582 49852 9588 49904
rect 9640 49852 9646 49904
rect 1762 49784 1768 49836
rect 1820 49784 1826 49836
rect 7098 49784 7104 49836
rect 7156 49824 7162 49836
rect 8021 49827 8079 49833
rect 8021 49824 8033 49827
rect 7156 49796 8033 49824
rect 7156 49784 7162 49796
rect 8021 49793 8033 49796
rect 8067 49793 8079 49827
rect 8021 49787 8079 49793
rect 9306 49784 9312 49836
rect 9364 49824 9370 49836
rect 9401 49827 9459 49833
rect 9401 49824 9413 49827
rect 9364 49796 9413 49824
rect 9364 49784 9370 49796
rect 9401 49793 9413 49796
rect 9447 49793 9459 49827
rect 9401 49787 9459 49793
rect 1670 49716 1676 49768
rect 1728 49756 1734 49768
rect 2225 49759 2283 49765
rect 2225 49756 2237 49759
rect 1728 49728 2237 49756
rect 1728 49716 1734 49728
rect 2225 49725 2237 49728
rect 2271 49725 2283 49759
rect 2225 49719 2283 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 1210 49240 1216 49292
rect 1268 49280 1274 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1268 49252 2053 49280
rect 1268 49240 1274 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 1578 49172 1584 49224
rect 1636 49172 1642 49224
rect 25038 49172 25044 49224
rect 25096 49172 25102 49224
rect 21450 49036 21456 49088
rect 21508 49076 21514 49088
rect 25225 49079 25283 49085
rect 25225 49076 25237 49079
rect 21508 49048 25237 49076
rect 21508 49036 21514 49048
rect 25225 49045 25237 49048
rect 25271 49045 25283 49079
rect 25225 49039 25283 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 11701 48875 11759 48881
rect 11701 48841 11713 48875
rect 11747 48872 11759 48875
rect 11974 48872 11980 48884
rect 11747 48844 11980 48872
rect 11747 48841 11759 48844
rect 11701 48835 11759 48841
rect 11974 48832 11980 48844
rect 12032 48832 12038 48884
rect 3970 48764 3976 48816
rect 4028 48804 4034 48816
rect 4249 48807 4307 48813
rect 4249 48804 4261 48807
rect 4028 48776 4261 48804
rect 4028 48764 4034 48776
rect 4249 48773 4261 48776
rect 4295 48773 4307 48807
rect 4249 48767 4307 48773
rect 3973 48671 4031 48677
rect 3973 48637 3985 48671
rect 4019 48637 4031 48671
rect 3973 48631 4031 48637
rect 3988 48532 4016 48631
rect 5368 48600 5396 48722
rect 11698 48696 11704 48748
rect 11756 48736 11762 48748
rect 11885 48739 11943 48745
rect 11885 48736 11897 48739
rect 11756 48708 11897 48736
rect 11756 48696 11762 48708
rect 11885 48705 11897 48708
rect 11931 48705 11943 48739
rect 11885 48699 11943 48705
rect 25038 48696 25044 48748
rect 25096 48696 25102 48748
rect 5997 48671 6055 48677
rect 5997 48637 6009 48671
rect 6043 48668 6055 48671
rect 9766 48668 9772 48680
rect 6043 48640 9772 48668
rect 6043 48637 6055 48640
rect 5997 48631 6055 48637
rect 9766 48628 9772 48640
rect 9824 48628 9830 48680
rect 10778 48600 10784 48612
rect 5368 48572 10784 48600
rect 10778 48560 10784 48572
rect 10836 48560 10842 48612
rect 9398 48532 9404 48544
rect 3988 48504 9404 48532
rect 9398 48492 9404 48504
rect 9456 48492 9462 48544
rect 25130 48492 25136 48544
rect 25188 48532 25194 48544
rect 25225 48535 25283 48541
rect 25225 48532 25237 48535
rect 25188 48504 25237 48532
rect 25188 48492 25194 48504
rect 25225 48501 25237 48504
rect 25271 48501 25283 48535
rect 25225 48495 25283 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 25038 48084 25044 48136
rect 25096 48084 25102 48136
rect 934 48016 940 48068
rect 992 48056 998 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 992 48028 1685 48056
rect 992 48016 998 48028
rect 1673 48025 1685 48028
rect 1719 48025 1731 48059
rect 1673 48019 1731 48025
rect 1857 48059 1915 48065
rect 1857 48025 1869 48059
rect 1903 48056 1915 48059
rect 3878 48056 3884 48068
rect 1903 48028 3884 48056
rect 1903 48025 1915 48028
rect 1857 48019 1915 48025
rect 3878 48016 3884 48028
rect 3936 48016 3942 48068
rect 25225 47991 25283 47997
rect 25225 47957 25237 47991
rect 25271 47988 25283 47991
rect 25406 47988 25412 48000
rect 25271 47960 25412 47988
rect 25271 47957 25283 47960
rect 25225 47951 25283 47957
rect 25406 47948 25412 47960
rect 25464 47948 25470 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 25038 47608 25044 47660
rect 25096 47608 25102 47660
rect 21358 47404 21364 47456
rect 21416 47444 21422 47456
rect 25225 47447 25283 47453
rect 25225 47444 25237 47447
rect 21416 47416 25237 47444
rect 21416 47404 21422 47416
rect 25225 47413 25237 47416
rect 25271 47413 25283 47447
rect 25225 47407 25283 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 6822 47200 6828 47252
rect 6880 47240 6886 47252
rect 9125 47243 9183 47249
rect 9125 47240 9137 47243
rect 6880 47212 9137 47240
rect 6880 47200 6886 47212
rect 9125 47209 9137 47212
rect 9171 47209 9183 47243
rect 9125 47203 9183 47209
rect 11517 47243 11575 47249
rect 11517 47209 11529 47243
rect 11563 47240 11575 47243
rect 11882 47240 11888 47252
rect 11563 47212 11888 47240
rect 11563 47209 11575 47212
rect 11517 47203 11575 47209
rect 11882 47200 11888 47212
rect 11940 47200 11946 47252
rect 15368 47243 15426 47249
rect 15368 47209 15380 47243
rect 15414 47240 15426 47243
rect 17402 47240 17408 47252
rect 15414 47212 17408 47240
rect 15414 47209 15426 47212
rect 15368 47203 15426 47209
rect 17402 47200 17408 47212
rect 17460 47200 17466 47252
rect 16390 47132 16396 47184
rect 16448 47172 16454 47184
rect 16448 47144 17908 47172
rect 16448 47132 16454 47144
rect 15105 47107 15163 47113
rect 15105 47073 15117 47107
rect 15151 47104 15163 47107
rect 15746 47104 15752 47116
rect 15151 47076 15752 47104
rect 15151 47073 15163 47076
rect 15105 47067 15163 47073
rect 15746 47064 15752 47076
rect 15804 47064 15810 47116
rect 16114 47064 16120 47116
rect 16172 47104 16178 47116
rect 17880 47113 17908 47144
rect 17865 47107 17923 47113
rect 16172 47076 17724 47104
rect 16172 47064 16178 47076
rect 9309 47039 9367 47045
rect 9309 47005 9321 47039
rect 9355 47036 9367 47039
rect 10594 47036 10600 47048
rect 9355 47008 10600 47036
rect 9355 47005 9367 47008
rect 9309 46999 9367 47005
rect 10594 46996 10600 47008
rect 10652 46996 10658 47048
rect 11606 46996 11612 47048
rect 11664 47036 11670 47048
rect 17696 47045 17724 47076
rect 17865 47073 17877 47107
rect 17911 47073 17923 47107
rect 17865 47067 17923 47073
rect 11701 47039 11759 47045
rect 11701 47036 11713 47039
rect 11664 47008 11713 47036
rect 11664 46996 11670 47008
rect 11701 47005 11713 47008
rect 11747 47005 11759 47039
rect 11701 46999 11759 47005
rect 17681 47039 17739 47045
rect 17681 47005 17693 47039
rect 17727 47005 17739 47039
rect 17681 46999 17739 47005
rect 15120 46940 15870 46968
rect 15010 46860 15016 46912
rect 15068 46900 15074 46912
rect 15120 46900 15148 46940
rect 16758 46928 16764 46980
rect 16816 46968 16822 46980
rect 16816 46940 16896 46968
rect 16816 46928 16822 46940
rect 16868 46909 16896 46940
rect 16942 46928 16948 46980
rect 17000 46968 17006 46980
rect 17770 46968 17776 46980
rect 17000 46940 17776 46968
rect 17000 46928 17006 46940
rect 17770 46928 17776 46940
rect 17828 46928 17834 46980
rect 15068 46872 15148 46900
rect 16853 46903 16911 46909
rect 15068 46860 15074 46872
rect 16853 46869 16865 46903
rect 16899 46869 16911 46903
rect 16853 46863 16911 46869
rect 17310 46860 17316 46912
rect 17368 46860 17374 46912
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7006 46656 7012 46708
rect 7064 46656 7070 46708
rect 15378 46656 15384 46708
rect 15436 46696 15442 46708
rect 16390 46696 16396 46708
rect 15436 46668 16396 46696
rect 15436 46656 15442 46668
rect 16390 46656 16396 46668
rect 16448 46656 16454 46708
rect 17218 46656 17224 46708
rect 17276 46656 17282 46708
rect 18509 46699 18567 46705
rect 18509 46665 18521 46699
rect 18555 46696 18567 46699
rect 18690 46696 18696 46708
rect 18555 46668 18696 46696
rect 18555 46665 18567 46668
rect 18509 46659 18567 46665
rect 18690 46656 18696 46668
rect 18748 46656 18754 46708
rect 17313 46631 17371 46637
rect 17313 46597 17325 46631
rect 17359 46628 17371 46631
rect 18874 46628 18880 46640
rect 17359 46600 18880 46628
rect 17359 46597 17371 46600
rect 17313 46591 17371 46597
rect 18524 46572 18552 46600
rect 18874 46588 18880 46600
rect 18932 46588 18938 46640
rect 7193 46563 7251 46569
rect 7193 46529 7205 46563
rect 7239 46560 7251 46563
rect 7834 46560 7840 46572
rect 7239 46532 7840 46560
rect 7239 46529 7251 46532
rect 7193 46523 7251 46529
rect 7834 46520 7840 46532
rect 7892 46520 7898 46572
rect 15010 46520 15016 46572
rect 15068 46520 15074 46572
rect 18414 46520 18420 46572
rect 18472 46520 18478 46572
rect 18506 46520 18512 46572
rect 18564 46520 18570 46572
rect 13354 46452 13360 46504
rect 13412 46492 13418 46504
rect 13633 46495 13691 46501
rect 13633 46492 13645 46495
rect 13412 46464 13645 46492
rect 13412 46452 13418 46464
rect 13633 46461 13645 46464
rect 13679 46461 13691 46495
rect 13633 46455 13691 46461
rect 13909 46495 13967 46501
rect 13909 46461 13921 46495
rect 13955 46492 13967 46495
rect 16022 46492 16028 46504
rect 13955 46464 16028 46492
rect 13955 46461 13967 46464
rect 13909 46455 13967 46461
rect 16022 46452 16028 46464
rect 16080 46452 16086 46504
rect 17402 46452 17408 46504
rect 17460 46452 17466 46504
rect 18690 46452 18696 46504
rect 18748 46452 18754 46504
rect 16853 46359 16911 46365
rect 16853 46325 16865 46359
rect 16899 46356 16911 46359
rect 17218 46356 17224 46368
rect 16899 46328 17224 46356
rect 16899 46325 16911 46328
rect 16853 46319 16911 46325
rect 17218 46316 17224 46328
rect 17276 46316 17282 46368
rect 17862 46316 17868 46368
rect 17920 46356 17926 46368
rect 18049 46359 18107 46365
rect 18049 46356 18061 46359
rect 17920 46328 18061 46356
rect 17920 46316 17926 46328
rect 18049 46325 18061 46328
rect 18095 46325 18107 46359
rect 18049 46319 18107 46325
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 5718 46112 5724 46164
rect 5776 46152 5782 46164
rect 7745 46155 7803 46161
rect 7745 46152 7757 46155
rect 5776 46124 7757 46152
rect 5776 46112 5782 46124
rect 7745 46121 7757 46124
rect 7791 46121 7803 46155
rect 7745 46115 7803 46121
rect 17402 46112 17408 46164
rect 17460 46152 17466 46164
rect 17589 46155 17647 46161
rect 17589 46152 17601 46155
rect 17460 46124 17601 46152
rect 17460 46112 17466 46124
rect 17589 46121 17601 46124
rect 17635 46121 17647 46155
rect 17589 46115 17647 46121
rect 20809 46087 20867 46093
rect 20809 46053 20821 46087
rect 20855 46084 20867 46087
rect 22462 46084 22468 46096
rect 20855 46056 22468 46084
rect 20855 46053 20867 46056
rect 20809 46047 20867 46053
rect 22462 46044 22468 46056
rect 22520 46044 22526 46096
rect 16117 46019 16175 46025
rect 16117 45985 16129 46019
rect 16163 46016 16175 46019
rect 17586 46016 17592 46028
rect 16163 45988 17592 46016
rect 16163 45985 16175 45988
rect 16117 45979 16175 45985
rect 17586 45976 17592 45988
rect 17644 45976 17650 46028
rect 19794 45976 19800 46028
rect 19852 46016 19858 46028
rect 19889 46019 19947 46025
rect 19889 46016 19901 46019
rect 19852 45988 19901 46016
rect 19852 45976 19858 45988
rect 19889 45985 19901 45988
rect 19935 45985 19947 46019
rect 19889 45979 19947 45985
rect 19978 45976 19984 46028
rect 20036 45976 20042 46028
rect 21453 46019 21511 46025
rect 21453 45985 21465 46019
rect 21499 46016 21511 46019
rect 22094 46016 22100 46028
rect 21499 45988 22100 46016
rect 21499 45985 21511 45988
rect 21453 45979 21511 45985
rect 22094 45976 22100 45988
rect 22152 45976 22158 46028
rect 934 45908 940 45960
rect 992 45948 998 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 992 45920 1593 45948
rect 992 45908 998 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 1857 45951 1915 45957
rect 1857 45917 1869 45951
rect 1903 45948 1915 45951
rect 9674 45948 9680 45960
rect 1903 45920 9680 45948
rect 1903 45917 1915 45920
rect 1857 45911 1915 45917
rect 9674 45908 9680 45920
rect 9732 45948 9738 45960
rect 9858 45948 9864 45960
rect 9732 45920 9864 45948
rect 9732 45908 9738 45920
rect 9858 45908 9864 45920
rect 9916 45908 9922 45960
rect 15838 45908 15844 45960
rect 15896 45908 15902 45960
rect 21269 45951 21327 45957
rect 21269 45917 21281 45951
rect 21315 45948 21327 45951
rect 22002 45948 22008 45960
rect 21315 45920 22008 45948
rect 21315 45917 21327 45920
rect 21269 45911 21327 45917
rect 22002 45908 22008 45920
rect 22060 45908 22066 45960
rect 24670 45908 24676 45960
rect 24728 45948 24734 45960
rect 25317 45951 25375 45957
rect 25317 45948 25329 45951
rect 24728 45920 25329 45948
rect 24728 45908 24734 45920
rect 25317 45917 25329 45920
rect 25363 45917 25375 45951
rect 25317 45911 25375 45917
rect 7282 45840 7288 45892
rect 7340 45880 7346 45892
rect 7653 45883 7711 45889
rect 7653 45880 7665 45883
rect 7340 45852 7665 45880
rect 7340 45840 7346 45852
rect 7653 45849 7665 45852
rect 7699 45849 7711 45883
rect 7653 45843 7711 45849
rect 16574 45840 16580 45892
rect 16632 45840 16638 45892
rect 19429 45815 19487 45821
rect 19429 45781 19441 45815
rect 19475 45812 19487 45815
rect 19610 45812 19616 45824
rect 19475 45784 19616 45812
rect 19475 45781 19487 45784
rect 19429 45775 19487 45781
rect 19610 45772 19616 45784
rect 19668 45772 19674 45824
rect 19794 45772 19800 45824
rect 19852 45772 19858 45824
rect 20622 45772 20628 45824
rect 20680 45812 20686 45824
rect 21177 45815 21235 45821
rect 21177 45812 21189 45815
rect 20680 45784 21189 45812
rect 20680 45772 20686 45784
rect 21177 45781 21189 45784
rect 21223 45781 21235 45815
rect 21177 45775 21235 45781
rect 22370 45772 22376 45824
rect 22428 45812 22434 45824
rect 25133 45815 25191 45821
rect 25133 45812 25145 45815
rect 22428 45784 25145 45812
rect 22428 45772 22434 45784
rect 25133 45781 25145 45784
rect 25179 45781 25191 45815
rect 25133 45775 25191 45781
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10965 45611 11023 45617
rect 10965 45577 10977 45611
rect 11011 45608 11023 45611
rect 11011 45580 11045 45608
rect 11011 45577 11023 45580
rect 10965 45571 11023 45577
rect 7190 45500 7196 45552
rect 7248 45540 7254 45552
rect 10980 45540 11008 45571
rect 15838 45568 15844 45620
rect 15896 45608 15902 45620
rect 15896 45580 16896 45608
rect 15896 45568 15902 45580
rect 13630 45540 13636 45552
rect 7248 45512 11008 45540
rect 11164 45512 13636 45540
rect 7248 45500 7254 45512
rect 7650 45432 7656 45484
rect 7708 45472 7714 45484
rect 8573 45475 8631 45481
rect 8573 45472 8585 45475
rect 7708 45444 8585 45472
rect 7708 45432 7714 45444
rect 8573 45441 8585 45444
rect 8619 45441 8631 45475
rect 8573 45435 8631 45441
rect 9953 45475 10011 45481
rect 9953 45441 9965 45475
rect 9999 45472 10011 45475
rect 10226 45472 10232 45484
rect 9999 45444 10232 45472
rect 9999 45441 10011 45444
rect 9953 45435 10011 45441
rect 10226 45432 10232 45444
rect 10284 45432 10290 45484
rect 11164 45481 11192 45512
rect 13630 45500 13636 45512
rect 13688 45500 13694 45552
rect 15010 45540 15016 45552
rect 14858 45512 15016 45540
rect 15010 45500 15016 45512
rect 15068 45500 15074 45552
rect 16868 45484 16896 45580
rect 18506 45540 18512 45552
rect 18354 45512 18512 45540
rect 18506 45500 18512 45512
rect 18564 45500 18570 45552
rect 19150 45500 19156 45552
rect 19208 45540 19214 45552
rect 20070 45540 20076 45552
rect 19208 45512 20076 45540
rect 19208 45500 19214 45512
rect 20070 45500 20076 45512
rect 20128 45500 20134 45552
rect 20165 45543 20223 45549
rect 20165 45509 20177 45543
rect 20211 45540 20223 45543
rect 21818 45540 21824 45552
rect 20211 45512 21824 45540
rect 20211 45509 20223 45512
rect 20165 45503 20223 45509
rect 21818 45500 21824 45512
rect 21876 45500 21882 45552
rect 11149 45475 11207 45481
rect 11149 45441 11161 45475
rect 11195 45441 11207 45475
rect 11149 45435 11207 45441
rect 11790 45432 11796 45484
rect 11848 45432 11854 45484
rect 16850 45432 16856 45484
rect 16908 45432 16914 45484
rect 24121 45475 24179 45481
rect 24121 45441 24133 45475
rect 24167 45472 24179 45475
rect 24578 45472 24584 45484
rect 24167 45444 24584 45472
rect 24167 45441 24179 45444
rect 24121 45435 24179 45441
rect 24578 45432 24584 45444
rect 24636 45432 24642 45484
rect 7466 45364 7472 45416
rect 7524 45404 7530 45416
rect 11977 45407 12035 45413
rect 11977 45404 11989 45407
rect 7524 45376 11989 45404
rect 7524 45364 7530 45376
rect 11977 45373 11989 45376
rect 12023 45373 12035 45407
rect 11977 45367 12035 45373
rect 13354 45364 13360 45416
rect 13412 45364 13418 45416
rect 13633 45407 13691 45413
rect 13633 45373 13645 45407
rect 13679 45404 13691 45407
rect 15378 45404 15384 45416
rect 13679 45376 15384 45404
rect 13679 45373 13691 45376
rect 13633 45367 13691 45373
rect 15378 45364 15384 45376
rect 15436 45364 15442 45416
rect 17129 45407 17187 45413
rect 17129 45373 17141 45407
rect 17175 45404 17187 45407
rect 18690 45404 18696 45416
rect 17175 45376 18696 45404
rect 17175 45373 17187 45376
rect 17129 45367 17187 45373
rect 18690 45364 18696 45376
rect 18748 45364 18754 45416
rect 20346 45364 20352 45416
rect 20404 45364 20410 45416
rect 24762 45364 24768 45416
rect 24820 45364 24826 45416
rect 8386 45296 8392 45348
rect 8444 45296 8450 45348
rect 9769 45339 9827 45345
rect 9769 45305 9781 45339
rect 9815 45336 9827 45339
rect 9950 45336 9956 45348
rect 9815 45308 9956 45336
rect 9815 45305 9827 45308
rect 9769 45299 9827 45305
rect 9950 45296 9956 45308
rect 10008 45296 10014 45348
rect 15102 45228 15108 45280
rect 15160 45228 15166 45280
rect 18598 45228 18604 45280
rect 18656 45228 18662 45280
rect 19702 45228 19708 45280
rect 19760 45228 19766 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 6362 45024 6368 45076
rect 6420 45064 6426 45076
rect 7561 45067 7619 45073
rect 7561 45064 7573 45067
rect 6420 45036 7573 45064
rect 6420 45024 6426 45036
rect 7561 45033 7573 45036
rect 7607 45033 7619 45067
rect 7561 45027 7619 45033
rect 9122 45024 9128 45076
rect 9180 45064 9186 45076
rect 10137 45067 10195 45073
rect 10137 45064 10149 45067
rect 9180 45036 10149 45064
rect 9180 45024 9186 45036
rect 10137 45033 10149 45036
rect 10183 45033 10195 45067
rect 10137 45027 10195 45033
rect 16022 45024 16028 45076
rect 16080 45064 16086 45076
rect 16390 45064 16396 45076
rect 16080 45036 16396 45064
rect 16080 45024 16086 45036
rect 16390 45024 16396 45036
rect 16448 45024 16454 45076
rect 24578 45024 24584 45076
rect 24636 45024 24642 45076
rect 21910 44888 21916 44940
rect 21968 44928 21974 44940
rect 22189 44931 22247 44937
rect 22189 44928 22201 44931
rect 21968 44900 22201 44928
rect 21968 44888 21974 44900
rect 22189 44897 22201 44900
rect 22235 44897 22247 44931
rect 22189 44891 22247 44897
rect 23290 44888 23296 44940
rect 23348 44888 23354 44940
rect 23474 44888 23480 44940
rect 23532 44888 23538 44940
rect 10686 44820 10692 44872
rect 10744 44820 10750 44872
rect 14274 44820 14280 44872
rect 14332 44820 14338 44872
rect 19426 44820 19432 44872
rect 19484 44820 19490 44872
rect 21266 44820 21272 44872
rect 21324 44860 21330 44872
rect 23201 44863 23259 44869
rect 23201 44860 23213 44863
rect 21324 44832 23213 44860
rect 21324 44820 21330 44832
rect 23201 44829 23213 44832
rect 23247 44829 23259 44863
rect 23201 44823 23259 44829
rect 23842 44820 23848 44872
rect 23900 44860 23906 44872
rect 24486 44860 24492 44872
rect 23900 44832 24492 44860
rect 23900 44820 23906 44832
rect 24486 44820 24492 44832
rect 24544 44860 24550 44872
rect 24765 44863 24823 44869
rect 24765 44860 24777 44863
rect 24544 44832 24777 44860
rect 24544 44820 24550 44832
rect 24765 44829 24777 44832
rect 24811 44829 24823 44863
rect 24765 44823 24823 44829
rect 7469 44795 7527 44801
rect 7469 44761 7481 44795
rect 7515 44792 7527 44795
rect 7558 44792 7564 44804
rect 7515 44764 7564 44792
rect 7515 44761 7527 44764
rect 7469 44755 7527 44761
rect 7558 44752 7564 44764
rect 7616 44752 7622 44804
rect 10045 44795 10103 44801
rect 10045 44761 10057 44795
rect 10091 44792 10103 44795
rect 10870 44792 10876 44804
rect 10091 44764 10876 44792
rect 10091 44761 10103 44764
rect 10045 44755 10103 44761
rect 10870 44752 10876 44764
rect 10928 44752 10934 44804
rect 10965 44795 11023 44801
rect 10965 44761 10977 44795
rect 11011 44792 11023 44795
rect 11054 44792 11060 44804
rect 11011 44764 11060 44792
rect 11011 44761 11023 44764
rect 10965 44755 11023 44761
rect 11054 44752 11060 44764
rect 11112 44752 11118 44804
rect 11348 44764 11454 44792
rect 9950 44684 9956 44736
rect 10008 44724 10014 44736
rect 10778 44724 10784 44736
rect 10008 44696 10784 44724
rect 10008 44684 10014 44696
rect 10778 44684 10784 44696
rect 10836 44724 10842 44736
rect 11348 44724 11376 44764
rect 14550 44752 14556 44804
rect 14608 44752 14614 44804
rect 15010 44792 15016 44804
rect 14660 44764 15016 44792
rect 10836 44696 11376 44724
rect 10836 44684 10842 44696
rect 12342 44684 12348 44736
rect 12400 44724 12406 44736
rect 12437 44727 12495 44733
rect 12437 44724 12449 44727
rect 12400 44696 12449 44724
rect 12400 44684 12406 44696
rect 12437 44693 12449 44696
rect 12483 44693 12495 44727
rect 12437 44687 12495 44693
rect 13814 44684 13820 44736
rect 13872 44724 13878 44736
rect 14660 44724 14688 44764
rect 15010 44752 15016 44764
rect 15068 44752 15074 44804
rect 19705 44795 19763 44801
rect 19705 44761 19717 44795
rect 19751 44792 19763 44795
rect 19794 44792 19800 44804
rect 19751 44764 19800 44792
rect 19751 44761 19763 44764
rect 19705 44755 19763 44761
rect 19794 44752 19800 44764
rect 19852 44792 19858 44804
rect 19978 44792 19984 44804
rect 19852 44764 19984 44792
rect 19852 44752 19858 44764
rect 19978 44752 19984 44764
rect 20036 44752 20042 44804
rect 20990 44792 20996 44804
rect 20930 44764 20996 44792
rect 20990 44752 20996 44764
rect 21048 44752 21054 44804
rect 21542 44752 21548 44804
rect 21600 44792 21606 44804
rect 22005 44795 22063 44801
rect 22005 44792 22017 44795
rect 21600 44764 22017 44792
rect 21600 44752 21606 44764
rect 22005 44761 22017 44764
rect 22051 44761 22063 44795
rect 22005 44755 22063 44761
rect 22097 44795 22155 44801
rect 22097 44761 22109 44795
rect 22143 44792 22155 44795
rect 23382 44792 23388 44804
rect 22143 44764 23388 44792
rect 22143 44761 22155 44764
rect 22097 44755 22155 44761
rect 23382 44752 23388 44764
rect 23440 44752 23446 44804
rect 13872 44696 14688 44724
rect 13872 44684 13878 44696
rect 19334 44684 19340 44736
rect 19392 44724 19398 44736
rect 21177 44727 21235 44733
rect 21177 44724 21189 44727
rect 19392 44696 21189 44724
rect 19392 44684 19398 44696
rect 21177 44693 21189 44696
rect 21223 44693 21235 44727
rect 21177 44687 21235 44693
rect 21634 44684 21640 44736
rect 21692 44684 21698 44736
rect 22830 44684 22836 44736
rect 22888 44684 22894 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 6270 44480 6276 44532
rect 6328 44520 6334 44532
rect 7285 44523 7343 44529
rect 7285 44520 7297 44523
rect 6328 44492 7297 44520
rect 6328 44480 6334 44492
rect 7285 44489 7297 44492
rect 7331 44489 7343 44523
rect 7285 44483 7343 44489
rect 8662 44480 8668 44532
rect 8720 44480 8726 44532
rect 11698 44480 11704 44532
rect 11756 44480 11762 44532
rect 12526 44480 12532 44532
rect 12584 44520 12590 44532
rect 14553 44523 14611 44529
rect 14553 44520 14565 44523
rect 12584 44492 14565 44520
rect 12584 44480 12590 44492
rect 14553 44489 14565 44492
rect 14599 44489 14611 44523
rect 14553 44483 14611 44489
rect 14645 44523 14703 44529
rect 14645 44489 14657 44523
rect 14691 44520 14703 44523
rect 15470 44520 15476 44532
rect 14691 44492 15476 44520
rect 14691 44489 14703 44492
rect 14645 44483 14703 44489
rect 15470 44480 15476 44492
rect 15528 44520 15534 44532
rect 16206 44520 16212 44532
rect 15528 44492 16212 44520
rect 15528 44480 15534 44492
rect 16206 44480 16212 44492
rect 16264 44480 16270 44532
rect 18690 44480 18696 44532
rect 18748 44520 18754 44532
rect 19429 44523 19487 44529
rect 19429 44520 19441 44523
rect 18748 44492 19441 44520
rect 18748 44480 18754 44492
rect 19429 44489 19441 44492
rect 19475 44489 19487 44523
rect 19429 44483 19487 44489
rect 20898 44480 20904 44532
rect 20956 44520 20962 44532
rect 21542 44520 21548 44532
rect 20956 44492 21548 44520
rect 20956 44480 20962 44492
rect 21542 44480 21548 44492
rect 21600 44480 21606 44532
rect 24489 44523 24547 44529
rect 24489 44520 24501 44523
rect 22066 44492 24501 44520
rect 9950 44412 9956 44464
rect 10008 44452 10014 44464
rect 10008 44424 10166 44452
rect 10008 44412 10014 44424
rect 18506 44412 18512 44464
rect 18564 44412 18570 44464
rect 22066 44452 22094 44492
rect 24489 44489 24501 44492
rect 24535 44489 24547 44523
rect 24489 44483 24547 44489
rect 23842 44452 23848 44464
rect 19720 44424 22094 44452
rect 23506 44424 23848 44452
rect 7190 44344 7196 44396
rect 7248 44344 7254 44396
rect 7742 44344 7748 44396
rect 7800 44384 7806 44396
rect 8021 44387 8079 44393
rect 8021 44384 8033 44387
rect 7800 44356 8033 44384
rect 7800 44344 7806 44356
rect 8021 44353 8033 44356
rect 8067 44353 8079 44387
rect 8021 44347 8079 44353
rect 8573 44387 8631 44393
rect 8573 44353 8585 44387
rect 8619 44384 8631 44387
rect 9030 44384 9036 44396
rect 8619 44356 9036 44384
rect 8619 44353 8631 44356
rect 8573 44347 8631 44353
rect 9030 44344 9036 44356
rect 9088 44344 9094 44396
rect 9398 44344 9404 44396
rect 9456 44344 9462 44396
rect 11974 44344 11980 44396
rect 12032 44384 12038 44396
rect 12069 44387 12127 44393
rect 12069 44384 12081 44387
rect 12032 44356 12081 44384
rect 12032 44344 12038 44356
rect 12069 44353 12081 44356
rect 12115 44353 12127 44387
rect 12069 44347 12127 44353
rect 12710 44344 12716 44396
rect 12768 44384 12774 44396
rect 12989 44387 13047 44393
rect 12989 44384 13001 44387
rect 12768 44356 13001 44384
rect 12768 44344 12774 44356
rect 12989 44353 13001 44356
rect 13035 44353 13047 44387
rect 12989 44347 13047 44353
rect 16850 44344 16856 44396
rect 16908 44384 16914 44396
rect 17681 44387 17739 44393
rect 17681 44384 17693 44387
rect 16908 44356 17693 44384
rect 16908 44344 16914 44356
rect 17681 44353 17693 44356
rect 17727 44353 17739 44387
rect 17681 44347 17739 44353
rect 9677 44319 9735 44325
rect 9677 44285 9689 44319
rect 9723 44316 9735 44319
rect 9766 44316 9772 44328
rect 9723 44288 9772 44316
rect 9723 44285 9735 44288
rect 9677 44279 9735 44285
rect 9766 44276 9772 44288
rect 9824 44316 9830 44328
rect 10042 44316 10048 44328
rect 9824 44288 10048 44316
rect 9824 44276 9830 44288
rect 10042 44276 10048 44288
rect 10100 44276 10106 44328
rect 10134 44276 10140 44328
rect 10192 44316 10198 44328
rect 10192 44288 10732 44316
rect 10192 44276 10198 44288
rect 6914 44208 6920 44260
rect 6972 44248 6978 44260
rect 7837 44251 7895 44257
rect 7837 44248 7849 44251
rect 6972 44220 7849 44248
rect 6972 44208 6978 44220
rect 7837 44217 7849 44220
rect 7883 44217 7895 44251
rect 10704 44248 10732 44288
rect 12158 44276 12164 44328
rect 12216 44276 12222 44328
rect 12342 44276 12348 44328
rect 12400 44276 12406 44328
rect 14829 44319 14887 44325
rect 14829 44285 14841 44319
rect 14875 44316 14887 44319
rect 14918 44316 14924 44328
rect 14875 44288 14924 44316
rect 14875 44285 14887 44288
rect 14829 44279 14887 44285
rect 14918 44276 14924 44288
rect 14976 44276 14982 44328
rect 17957 44319 18015 44325
rect 17957 44285 17969 44319
rect 18003 44316 18015 44319
rect 19518 44316 19524 44328
rect 18003 44288 19524 44316
rect 18003 44285 18015 44288
rect 17957 44279 18015 44285
rect 19518 44276 19524 44288
rect 19576 44276 19582 44328
rect 13173 44251 13231 44257
rect 13173 44248 13185 44251
rect 10704 44220 13185 44248
rect 7837 44211 7895 44217
rect 13173 44217 13185 44220
rect 13219 44217 13231 44251
rect 13173 44211 13231 44217
rect 9766 44140 9772 44192
rect 9824 44180 9830 44192
rect 10226 44180 10232 44192
rect 9824 44152 10232 44180
rect 9824 44140 9830 44152
rect 10226 44140 10232 44152
rect 10284 44140 10290 44192
rect 11054 44140 11060 44192
rect 11112 44180 11118 44192
rect 11149 44183 11207 44189
rect 11149 44180 11161 44183
rect 11112 44152 11161 44180
rect 11112 44140 11118 44152
rect 11149 44149 11161 44152
rect 11195 44180 11207 44183
rect 12250 44180 12256 44192
rect 11195 44152 12256 44180
rect 11195 44149 11207 44152
rect 11149 44143 11207 44149
rect 12250 44140 12256 44152
rect 12308 44140 12314 44192
rect 14182 44140 14188 44192
rect 14240 44140 14246 44192
rect 14550 44140 14556 44192
rect 14608 44180 14614 44192
rect 16758 44180 16764 44192
rect 14608 44152 16764 44180
rect 14608 44140 14614 44152
rect 16758 44140 16764 44152
rect 16816 44180 16822 44192
rect 17402 44180 17408 44192
rect 16816 44152 17408 44180
rect 16816 44140 16822 44152
rect 17402 44140 17408 44152
rect 17460 44140 17466 44192
rect 18414 44140 18420 44192
rect 18472 44180 18478 44192
rect 19720 44180 19748 44424
rect 23842 44412 23848 44424
rect 23900 44412 23906 44464
rect 24673 44387 24731 44393
rect 24673 44353 24685 44387
rect 24719 44384 24731 44387
rect 24854 44384 24860 44396
rect 24719 44356 24860 44384
rect 24719 44353 24731 44356
rect 24673 44347 24731 44353
rect 24854 44344 24860 44356
rect 24912 44344 24918 44396
rect 25314 44344 25320 44396
rect 25372 44344 25378 44396
rect 22002 44276 22008 44328
rect 22060 44276 22066 44328
rect 22278 44276 22284 44328
rect 22336 44276 22342 44328
rect 18472 44152 19748 44180
rect 18472 44140 18478 44152
rect 20346 44140 20352 44192
rect 20404 44180 20410 44192
rect 23753 44183 23811 44189
rect 23753 44180 23765 44183
rect 20404 44152 23765 44180
rect 20404 44140 20410 44152
rect 23753 44149 23765 44152
rect 23799 44149 23811 44183
rect 23753 44143 23811 44149
rect 24946 44140 24952 44192
rect 25004 44180 25010 44192
rect 25133 44183 25191 44189
rect 25133 44180 25145 44183
rect 25004 44152 25145 44180
rect 25004 44140 25010 44152
rect 25133 44149 25145 44152
rect 25179 44149 25191 44183
rect 25133 44143 25191 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 6546 43936 6552 43988
rect 6604 43936 6610 43988
rect 7374 43936 7380 43988
rect 7432 43976 7438 43988
rect 8481 43979 8539 43985
rect 8481 43976 8493 43979
rect 7432 43948 8493 43976
rect 7432 43936 7438 43948
rect 8481 43945 8493 43948
rect 8527 43945 8539 43979
rect 8481 43939 8539 43945
rect 8938 43936 8944 43988
rect 8996 43976 9002 43988
rect 9861 43979 9919 43985
rect 9861 43976 9873 43979
rect 8996 43948 9873 43976
rect 8996 43936 9002 43948
rect 9861 43945 9873 43948
rect 9907 43945 9919 43979
rect 9861 43939 9919 43945
rect 17586 43936 17592 43988
rect 17644 43936 17650 43988
rect 19794 43936 19800 43988
rect 19852 43976 19858 43988
rect 21177 43979 21235 43985
rect 21177 43976 21189 43979
rect 19852 43948 21189 43976
rect 19852 43936 19858 43948
rect 21177 43945 21189 43948
rect 21223 43945 21235 43979
rect 21177 43939 21235 43945
rect 9214 43868 9220 43920
rect 9272 43908 9278 43920
rect 10689 43911 10747 43917
rect 10689 43908 10701 43911
rect 9272 43880 10701 43908
rect 9272 43868 9278 43880
rect 10689 43877 10701 43880
rect 10735 43877 10747 43911
rect 10689 43871 10747 43877
rect 16117 43843 16175 43849
rect 16117 43809 16129 43843
rect 16163 43840 16175 43843
rect 16206 43840 16212 43852
rect 16163 43812 16212 43840
rect 16163 43809 16175 43812
rect 16117 43803 16175 43809
rect 16206 43800 16212 43812
rect 16264 43840 16270 43852
rect 18598 43840 18604 43852
rect 16264 43812 18604 43840
rect 16264 43800 16270 43812
rect 18598 43800 18604 43812
rect 18656 43800 18662 43852
rect 19705 43843 19763 43849
rect 19705 43809 19717 43843
rect 19751 43840 19763 43843
rect 20070 43840 20076 43852
rect 19751 43812 20076 43840
rect 19751 43809 19763 43812
rect 19705 43803 19763 43809
rect 20070 43800 20076 43812
rect 20128 43800 20134 43852
rect 25130 43840 25136 43852
rect 21100 43812 25136 43840
rect 8389 43775 8447 43781
rect 8389 43741 8401 43775
rect 8435 43772 8447 43775
rect 10318 43772 10324 43784
rect 8435 43744 10324 43772
rect 8435 43741 8447 43744
rect 8389 43735 8447 43741
rect 10318 43732 10324 43744
rect 10376 43732 10382 43784
rect 10686 43732 10692 43784
rect 10744 43772 10750 43784
rect 11790 43772 11796 43784
rect 10744 43744 11796 43772
rect 10744 43732 10750 43744
rect 11790 43732 11796 43744
rect 11848 43732 11854 43784
rect 13814 43772 13820 43784
rect 13202 43758 13820 43772
rect 13188 43744 13820 43758
rect 6457 43707 6515 43713
rect 6457 43673 6469 43707
rect 6503 43704 6515 43707
rect 8294 43704 8300 43716
rect 6503 43676 8300 43704
rect 6503 43673 6515 43676
rect 6457 43667 6515 43673
rect 8294 43664 8300 43676
rect 8352 43664 8358 43716
rect 9769 43707 9827 43713
rect 9769 43673 9781 43707
rect 9815 43704 9827 43707
rect 10226 43704 10232 43716
rect 9815 43676 10232 43704
rect 9815 43673 9827 43676
rect 9769 43667 9827 43673
rect 10226 43664 10232 43676
rect 10284 43664 10290 43716
rect 10502 43664 10508 43716
rect 10560 43664 10566 43716
rect 12069 43707 12127 43713
rect 12069 43673 12081 43707
rect 12115 43704 12127 43707
rect 12342 43704 12348 43716
rect 12115 43676 12348 43704
rect 12115 43673 12127 43676
rect 12069 43667 12127 43673
rect 12342 43664 12348 43676
rect 12400 43664 12406 43716
rect 9950 43596 9956 43648
rect 10008 43636 10014 43648
rect 13188 43636 13216 43744
rect 13814 43732 13820 43744
rect 13872 43732 13878 43784
rect 15286 43732 15292 43784
rect 15344 43772 15350 43784
rect 15838 43772 15844 43784
rect 15344 43744 15844 43772
rect 15344 43732 15350 43744
rect 15838 43732 15844 43744
rect 15896 43732 15902 43784
rect 18782 43732 18788 43784
rect 18840 43772 18846 43784
rect 19429 43775 19487 43781
rect 19429 43772 19441 43775
rect 18840 43744 19441 43772
rect 18840 43732 18846 43744
rect 19429 43741 19441 43744
rect 19475 43741 19487 43775
rect 19429 43735 19487 43741
rect 16574 43664 16580 43716
rect 16632 43664 16638 43716
rect 20990 43704 20996 43716
rect 20930 43676 20996 43704
rect 20990 43664 20996 43676
rect 21048 43664 21054 43716
rect 10008 43608 13216 43636
rect 10008 43596 10014 43608
rect 13538 43596 13544 43648
rect 13596 43596 13602 43648
rect 17494 43596 17500 43648
rect 17552 43636 17558 43648
rect 21100 43636 21128 43812
rect 25130 43800 25136 43812
rect 25188 43800 25194 43852
rect 22002 43732 22008 43784
rect 22060 43772 22066 43784
rect 22189 43775 22247 43781
rect 22189 43772 22201 43775
rect 22060 43744 22201 43772
rect 22060 43732 22066 43744
rect 22189 43741 22201 43744
rect 22235 43741 22247 43775
rect 22189 43735 22247 43741
rect 24762 43732 24768 43784
rect 24820 43772 24826 43784
rect 25317 43775 25375 43781
rect 25317 43772 25329 43775
rect 24820 43744 25329 43772
rect 24820 43732 24826 43744
rect 25317 43741 25329 43744
rect 25363 43741 25375 43775
rect 25317 43735 25375 43741
rect 22465 43707 22523 43713
rect 22465 43704 22477 43707
rect 22204 43676 22477 43704
rect 22204 43648 22232 43676
rect 22465 43673 22477 43676
rect 22511 43673 22523 43707
rect 23842 43704 23848 43716
rect 23690 43676 23848 43704
rect 22465 43667 22523 43673
rect 23842 43664 23848 43676
rect 23900 43664 23906 43716
rect 17552 43608 21128 43636
rect 17552 43596 17558 43608
rect 22186 43596 22192 43648
rect 22244 43596 22250 43648
rect 22278 43596 22284 43648
rect 22336 43636 22342 43648
rect 23937 43639 23995 43645
rect 23937 43636 23949 43639
rect 22336 43608 23949 43636
rect 22336 43596 22342 43608
rect 23937 43605 23949 43608
rect 23983 43605 23995 43639
rect 23937 43599 23995 43605
rect 25133 43639 25191 43645
rect 25133 43605 25145 43639
rect 25179 43636 25191 43639
rect 25498 43636 25504 43648
rect 25179 43608 25504 43636
rect 25179 43605 25191 43608
rect 25133 43599 25191 43605
rect 25498 43596 25504 43608
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 5534 43392 5540 43444
rect 5592 43392 5598 43444
rect 10686 43432 10692 43444
rect 8588 43404 10692 43432
rect 5166 43256 5172 43308
rect 5224 43296 5230 43308
rect 8588 43305 8616 43404
rect 10686 43392 10692 43404
rect 10744 43392 10750 43444
rect 12158 43392 12164 43444
rect 12216 43432 12222 43444
rect 12253 43435 12311 43441
rect 12253 43432 12265 43435
rect 12216 43404 12265 43432
rect 12216 43392 12222 43404
rect 12253 43401 12265 43404
rect 12299 43401 12311 43435
rect 12253 43395 12311 43401
rect 17218 43392 17224 43444
rect 17276 43432 17282 43444
rect 17313 43435 17371 43441
rect 17313 43432 17325 43435
rect 17276 43404 17325 43432
rect 17276 43392 17282 43404
rect 17313 43401 17325 43404
rect 17359 43401 17371 43435
rect 17313 43395 17371 43401
rect 22186 43392 22192 43444
rect 22244 43432 22250 43444
rect 23753 43435 23811 43441
rect 23753 43432 23765 43435
rect 22244 43404 23765 43432
rect 22244 43392 22250 43404
rect 23753 43401 23765 43404
rect 23799 43401 23811 43435
rect 23753 43395 23811 43401
rect 9490 43324 9496 43376
rect 9548 43324 9554 43376
rect 23842 43364 23848 43376
rect 23506 43336 23848 43364
rect 23842 43324 23848 43336
rect 23900 43324 23906 43376
rect 5721 43299 5779 43305
rect 5721 43296 5733 43299
rect 5224 43268 5733 43296
rect 5224 43256 5230 43268
rect 5721 43265 5733 43268
rect 5767 43265 5779 43299
rect 5721 43259 5779 43265
rect 8573 43299 8631 43305
rect 8573 43265 8585 43299
rect 8619 43265 8631 43299
rect 8573 43259 8631 43265
rect 12621 43299 12679 43305
rect 12621 43265 12633 43299
rect 12667 43296 12679 43299
rect 15194 43296 15200 43308
rect 12667 43268 15200 43296
rect 12667 43265 12679 43268
rect 12621 43259 12679 43265
rect 15194 43256 15200 43268
rect 15252 43256 15258 43308
rect 17221 43299 17279 43305
rect 17221 43265 17233 43299
rect 17267 43296 17279 43299
rect 17494 43296 17500 43308
rect 17267 43268 17500 43296
rect 17267 43265 17279 43268
rect 17221 43259 17279 43265
rect 17494 43256 17500 43268
rect 17552 43296 17558 43308
rect 17678 43296 17684 43308
rect 17552 43268 17684 43296
rect 17552 43256 17558 43268
rect 17678 43256 17684 43268
rect 17736 43256 17742 43308
rect 24489 43299 24547 43305
rect 24489 43265 24501 43299
rect 24535 43296 24547 43299
rect 24854 43296 24860 43308
rect 24535 43268 24860 43296
rect 24535 43265 24547 43268
rect 24489 43259 24547 43265
rect 24854 43256 24860 43268
rect 24912 43256 24918 43308
rect 8849 43231 8907 43237
rect 8849 43197 8861 43231
rect 8895 43228 8907 43231
rect 8895 43200 9996 43228
rect 8895 43197 8907 43200
rect 8849 43191 8907 43197
rect 9968 43160 9996 43200
rect 10042 43188 10048 43240
rect 10100 43228 10106 43240
rect 12713 43231 12771 43237
rect 12713 43228 12725 43231
rect 10100 43200 12725 43228
rect 10100 43188 10106 43200
rect 12713 43197 12725 43200
rect 12759 43197 12771 43231
rect 12713 43191 12771 43197
rect 12805 43231 12863 43237
rect 12805 43197 12817 43231
rect 12851 43197 12863 43231
rect 12805 43191 12863 43197
rect 9968 43132 12296 43160
rect 9490 43052 9496 43104
rect 9548 43092 9554 43104
rect 9950 43092 9956 43104
rect 9548 43064 9956 43092
rect 9548 43052 9554 43064
rect 9950 43052 9956 43064
rect 10008 43052 10014 43104
rect 10321 43095 10379 43101
rect 10321 43061 10333 43095
rect 10367 43092 10379 43095
rect 10410 43092 10416 43104
rect 10367 43064 10416 43092
rect 10367 43061 10379 43064
rect 10321 43055 10379 43061
rect 10410 43052 10416 43064
rect 10468 43052 10474 43104
rect 12268 43092 12296 43132
rect 12342 43120 12348 43172
rect 12400 43160 12406 43172
rect 12820 43160 12848 43191
rect 17402 43188 17408 43240
rect 17460 43188 17466 43240
rect 22002 43188 22008 43240
rect 22060 43188 22066 43240
rect 22281 43231 22339 43237
rect 22281 43228 22293 43231
rect 22112 43200 22293 43228
rect 12400 43132 12848 43160
rect 12400 43120 12406 43132
rect 22112 43104 22140 43200
rect 22281 43197 22293 43200
rect 22327 43228 22339 43231
rect 22646 43228 22652 43240
rect 22327 43200 22652 43228
rect 22327 43197 22339 43200
rect 22281 43191 22339 43197
rect 22646 43188 22652 43200
rect 22704 43188 22710 43240
rect 23750 43188 23756 43240
rect 23808 43228 23814 43240
rect 24765 43231 24823 43237
rect 24765 43228 24777 43231
rect 23808 43200 24777 43228
rect 23808 43188 23814 43200
rect 24765 43197 24777 43200
rect 24811 43197 24823 43231
rect 24765 43191 24823 43197
rect 15378 43092 15384 43104
rect 12268 43064 15384 43092
rect 15378 43052 15384 43064
rect 15436 43052 15442 43104
rect 16666 43052 16672 43104
rect 16724 43092 16730 43104
rect 16853 43095 16911 43101
rect 16853 43092 16865 43095
rect 16724 43064 16865 43092
rect 16724 43052 16730 43064
rect 16853 43061 16865 43064
rect 16899 43061 16911 43095
rect 16853 43055 16911 43061
rect 22094 43052 22100 43104
rect 22152 43052 22158 43104
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 13814 42848 13820 42900
rect 13872 42888 13878 42900
rect 14540 42891 14598 42897
rect 14540 42888 14552 42891
rect 13872 42860 14552 42888
rect 13872 42848 13878 42860
rect 14540 42857 14552 42860
rect 14586 42888 14598 42891
rect 15102 42888 15108 42900
rect 14586 42860 15108 42888
rect 14586 42857 14598 42860
rect 14540 42851 14598 42857
rect 15102 42848 15108 42860
rect 15160 42848 15166 42900
rect 19692 42891 19750 42897
rect 19692 42857 19704 42891
rect 19738 42888 19750 42891
rect 20346 42888 20352 42900
rect 19738 42860 20352 42888
rect 19738 42857 19750 42860
rect 19692 42851 19750 42857
rect 20346 42848 20352 42860
rect 20404 42848 20410 42900
rect 20990 42848 20996 42900
rect 21048 42888 21054 42900
rect 23842 42888 23848 42900
rect 21048 42860 23848 42888
rect 21048 42848 21054 42860
rect 23842 42848 23848 42860
rect 23900 42848 23906 42900
rect 10226 42820 10232 42832
rect 10060 42792 10232 42820
rect 3694 42712 3700 42764
rect 3752 42752 3758 42764
rect 4433 42755 4491 42761
rect 4433 42752 4445 42755
rect 3752 42724 4445 42752
rect 3752 42712 3758 42724
rect 4433 42721 4445 42724
rect 4479 42721 4491 42755
rect 4433 42715 4491 42721
rect 6454 42712 6460 42764
rect 6512 42752 6518 42764
rect 10060 42761 10088 42792
rect 10226 42780 10232 42792
rect 10284 42780 10290 42832
rect 18598 42820 18604 42832
rect 18156 42792 18604 42820
rect 6549 42755 6607 42761
rect 6549 42752 6561 42755
rect 6512 42724 6561 42752
rect 6512 42712 6518 42724
rect 6549 42721 6561 42724
rect 6595 42721 6607 42755
rect 8573 42755 8631 42761
rect 8573 42752 8585 42755
rect 6549 42715 6607 42721
rect 6886 42724 8585 42752
rect 5350 42644 5356 42696
rect 5408 42684 5414 42696
rect 6886 42684 6914 42724
rect 8573 42721 8585 42724
rect 8619 42721 8631 42755
rect 8573 42715 8631 42721
rect 10045 42755 10103 42761
rect 10045 42721 10057 42755
rect 10091 42721 10103 42755
rect 10045 42715 10103 42721
rect 12618 42712 12624 42764
rect 12676 42712 12682 42764
rect 14274 42712 14280 42764
rect 14332 42712 14338 42764
rect 17862 42712 17868 42764
rect 17920 42752 17926 42764
rect 18156 42761 18184 42792
rect 18598 42780 18604 42792
rect 18656 42780 18662 42832
rect 17957 42755 18015 42761
rect 17957 42752 17969 42755
rect 17920 42724 17969 42752
rect 17920 42712 17926 42724
rect 17957 42721 17969 42724
rect 18003 42721 18015 42755
rect 17957 42715 18015 42721
rect 18141 42755 18199 42761
rect 18141 42721 18153 42755
rect 18187 42721 18199 42755
rect 18141 42715 18199 42721
rect 19426 42712 19432 42764
rect 19484 42752 19490 42764
rect 21266 42752 21272 42764
rect 19484 42724 21272 42752
rect 19484 42712 19490 42724
rect 21266 42712 21272 42724
rect 21324 42752 21330 42764
rect 22002 42752 22008 42764
rect 21324 42724 22008 42752
rect 21324 42712 21330 42724
rect 22002 42712 22008 42724
rect 22060 42752 22066 42764
rect 22281 42755 22339 42761
rect 22281 42752 22293 42755
rect 22060 42724 22293 42752
rect 22060 42712 22066 42724
rect 22281 42721 22293 42724
rect 22327 42721 22339 42755
rect 22281 42715 22339 42721
rect 5408 42656 6914 42684
rect 5408 42644 5414 42656
rect 7098 42644 7104 42696
rect 7156 42684 7162 42696
rect 7193 42687 7251 42693
rect 7193 42684 7205 42687
rect 7156 42656 7205 42684
rect 7156 42644 7162 42656
rect 7193 42653 7205 42656
rect 7239 42653 7251 42687
rect 7193 42647 7251 42653
rect 7837 42687 7895 42693
rect 7837 42653 7849 42687
rect 7883 42653 7895 42687
rect 7837 42647 7895 42653
rect 9769 42687 9827 42693
rect 9769 42653 9781 42687
rect 9815 42684 9827 42687
rect 9858 42684 9864 42696
rect 9815 42656 9864 42684
rect 9815 42653 9827 42656
rect 9769 42647 9827 42653
rect 4154 42576 4160 42628
rect 4212 42616 4218 42628
rect 4249 42619 4307 42625
rect 4249 42616 4261 42619
rect 4212 42588 4261 42616
rect 4212 42576 4218 42588
rect 4249 42585 4261 42588
rect 4295 42585 4307 42619
rect 4249 42579 4307 42585
rect 6365 42619 6423 42625
rect 6365 42585 6377 42619
rect 6411 42616 6423 42619
rect 6454 42616 6460 42628
rect 6411 42588 6460 42616
rect 6411 42585 6423 42588
rect 6365 42579 6423 42585
rect 6454 42576 6460 42588
rect 6512 42576 6518 42628
rect 6914 42576 6920 42628
rect 6972 42616 6978 42628
rect 7852 42616 7880 42647
rect 9858 42644 9864 42656
rect 9916 42644 9922 42696
rect 11790 42644 11796 42696
rect 11848 42684 11854 42696
rect 14292 42684 14320 42712
rect 11848 42656 14320 42684
rect 11848 42644 11854 42656
rect 25314 42644 25320 42696
rect 25372 42644 25378 42696
rect 6972 42588 7880 42616
rect 8389 42619 8447 42625
rect 6972 42576 6978 42588
rect 8389 42585 8401 42619
rect 8435 42616 8447 42619
rect 8570 42616 8576 42628
rect 8435 42588 8576 42616
rect 8435 42585 8447 42588
rect 8389 42579 8447 42585
rect 8570 42576 8576 42588
rect 8628 42576 8634 42628
rect 10042 42616 10048 42628
rect 9416 42588 10048 42616
rect 7006 42508 7012 42560
rect 7064 42508 7070 42560
rect 7653 42551 7711 42557
rect 7653 42517 7665 42551
rect 7699 42548 7711 42551
rect 9306 42548 9312 42560
rect 7699 42520 9312 42548
rect 7699 42517 7711 42520
rect 7653 42511 7711 42517
rect 9306 42508 9312 42520
rect 9364 42508 9370 42560
rect 9416 42557 9444 42588
rect 10042 42576 10048 42588
rect 10100 42576 10106 42628
rect 11514 42576 11520 42628
rect 11572 42616 11578 42628
rect 12345 42619 12403 42625
rect 12345 42616 12357 42619
rect 11572 42588 12357 42616
rect 11572 42576 11578 42588
rect 12345 42585 12357 42588
rect 12391 42585 12403 42619
rect 12345 42579 12403 42585
rect 14274 42576 14280 42628
rect 14332 42616 14338 42628
rect 16758 42616 16764 42628
rect 14332 42588 15042 42616
rect 15948 42588 16764 42616
rect 14332 42576 14338 42588
rect 9401 42551 9459 42557
rect 9401 42517 9413 42551
rect 9447 42517 9459 42551
rect 9401 42511 9459 42517
rect 9861 42551 9919 42557
rect 9861 42517 9873 42551
rect 9907 42548 9919 42551
rect 9950 42548 9956 42560
rect 9907 42520 9956 42548
rect 9907 42517 9919 42520
rect 9861 42511 9919 42517
rect 9950 42508 9956 42520
rect 10008 42548 10014 42560
rect 10134 42548 10140 42560
rect 10008 42520 10140 42548
rect 10008 42508 10014 42520
rect 10134 42508 10140 42520
rect 10192 42508 10198 42560
rect 10594 42508 10600 42560
rect 10652 42548 10658 42560
rect 11977 42551 12035 42557
rect 11977 42548 11989 42551
rect 10652 42520 11989 42548
rect 10652 42508 10658 42520
rect 11977 42517 11989 42520
rect 12023 42517 12035 42551
rect 11977 42511 12035 42517
rect 12437 42551 12495 42557
rect 12437 42517 12449 42551
rect 12483 42548 12495 42551
rect 15948 42548 15976 42588
rect 16758 42576 16764 42588
rect 16816 42576 16822 42628
rect 20990 42616 20996 42628
rect 20930 42588 20996 42616
rect 20990 42576 20996 42588
rect 21048 42576 21054 42628
rect 22554 42576 22560 42628
rect 22612 42576 22618 42628
rect 23842 42616 23848 42628
rect 23782 42588 23848 42616
rect 23842 42576 23848 42588
rect 23900 42616 23906 42628
rect 24578 42616 24584 42628
rect 23900 42588 24584 42616
rect 23900 42576 23906 42588
rect 24578 42576 24584 42588
rect 24636 42576 24642 42628
rect 12483 42520 15976 42548
rect 12483 42517 12495 42520
rect 12437 42511 12495 42517
rect 16022 42508 16028 42560
rect 16080 42508 16086 42560
rect 17494 42508 17500 42560
rect 17552 42508 17558 42560
rect 17770 42508 17776 42560
rect 17828 42548 17834 42560
rect 17865 42551 17923 42557
rect 17865 42548 17877 42551
rect 17828 42520 17877 42548
rect 17828 42508 17834 42520
rect 17865 42517 17877 42520
rect 17911 42517 17923 42551
rect 17865 42511 17923 42517
rect 21174 42508 21180 42560
rect 21232 42508 21238 42560
rect 23566 42508 23572 42560
rect 23624 42548 23630 42560
rect 24029 42551 24087 42557
rect 24029 42548 24041 42551
rect 23624 42520 24041 42548
rect 23624 42508 23630 42520
rect 24029 42517 24041 42520
rect 24075 42517 24087 42551
rect 24029 42511 24087 42517
rect 25133 42551 25191 42557
rect 25133 42517 25145 42551
rect 25179 42548 25191 42551
rect 25222 42548 25228 42560
rect 25179 42520 25228 42548
rect 25179 42517 25191 42520
rect 25133 42511 25191 42517
rect 25222 42508 25228 42520
rect 25280 42508 25286 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 1762 42304 1768 42356
rect 1820 42344 1826 42356
rect 3881 42347 3939 42353
rect 3881 42344 3893 42347
rect 1820 42316 3893 42344
rect 1820 42304 1826 42316
rect 3881 42313 3893 42316
rect 3927 42313 3939 42347
rect 9490 42344 9496 42356
rect 3881 42307 3939 42313
rect 8496 42316 9496 42344
rect 8386 42236 8392 42288
rect 8444 42276 8450 42288
rect 8496 42276 8524 42316
rect 9490 42304 9496 42316
rect 9548 42304 9554 42356
rect 11606 42304 11612 42356
rect 11664 42344 11670 42356
rect 11701 42347 11759 42353
rect 11701 42344 11713 42347
rect 11664 42316 11713 42344
rect 11664 42304 11670 42316
rect 11701 42313 11713 42316
rect 11747 42313 11759 42347
rect 11701 42307 11759 42313
rect 19518 42304 19524 42356
rect 19576 42344 19582 42356
rect 19613 42347 19671 42353
rect 19613 42344 19625 42347
rect 19576 42316 19625 42344
rect 19576 42304 19582 42316
rect 19613 42313 19625 42316
rect 19659 42344 19671 42347
rect 20438 42344 20444 42356
rect 19659 42316 20444 42344
rect 19659 42313 19671 42316
rect 19613 42307 19671 42313
rect 20438 42304 20444 42316
rect 20496 42304 20502 42356
rect 22462 42304 22468 42356
rect 22520 42304 22526 42356
rect 12161 42279 12219 42285
rect 8444 42248 8602 42276
rect 8444 42236 8450 42248
rect 12161 42245 12173 42279
rect 12207 42276 12219 42279
rect 12250 42276 12256 42288
rect 12207 42248 12256 42276
rect 12207 42245 12219 42248
rect 12161 42239 12219 42245
rect 12250 42236 12256 42248
rect 12308 42236 12314 42288
rect 14366 42236 14372 42288
rect 14424 42236 14430 42288
rect 18598 42236 18604 42288
rect 18656 42236 18662 42288
rect 21266 42236 21272 42288
rect 21324 42276 21330 42288
rect 22002 42276 22008 42288
rect 21324 42248 22008 42276
rect 21324 42236 21330 42248
rect 22002 42236 22008 42248
rect 22060 42276 22066 42288
rect 22060 42248 23336 42276
rect 22060 42236 22066 42248
rect 3786 42168 3792 42220
rect 3844 42168 3850 42220
rect 11882 42168 11888 42220
rect 11940 42208 11946 42220
rect 12069 42211 12127 42217
rect 12069 42208 12081 42211
rect 11940 42180 12081 42208
rect 11940 42168 11946 42180
rect 12069 42177 12081 42180
rect 12115 42177 12127 42211
rect 12069 42171 12127 42177
rect 15286 42168 15292 42220
rect 15344 42208 15350 42220
rect 17862 42208 17868 42220
rect 15344 42180 17868 42208
rect 15344 42168 15350 42180
rect 17862 42168 17868 42180
rect 17920 42168 17926 42220
rect 19426 42168 19432 42220
rect 19484 42208 19490 42220
rect 20533 42211 20591 42217
rect 20533 42208 20545 42211
rect 19484 42180 20545 42208
rect 19484 42168 19490 42180
rect 20533 42177 20545 42180
rect 20579 42177 20591 42211
rect 20533 42171 20591 42177
rect 20714 42168 20720 42220
rect 20772 42208 20778 42220
rect 23308 42217 23336 42248
rect 23566 42236 23572 42288
rect 23624 42236 23630 42288
rect 24578 42236 24584 42288
rect 24636 42236 24642 42288
rect 22373 42211 22431 42217
rect 22373 42208 22385 42211
rect 20772 42180 22385 42208
rect 20772 42168 20778 42180
rect 22373 42177 22385 42180
rect 22419 42177 22431 42211
rect 22373 42171 22431 42177
rect 23293 42211 23351 42217
rect 23293 42177 23305 42211
rect 23339 42177 23351 42211
rect 23293 42171 23351 42177
rect 7837 42143 7895 42149
rect 7837 42109 7849 42143
rect 7883 42109 7895 42143
rect 7837 42103 7895 42109
rect 8113 42143 8171 42149
rect 8113 42109 8125 42143
rect 8159 42140 8171 42143
rect 8478 42140 8484 42152
rect 8159 42112 8484 42140
rect 8159 42109 8171 42112
rect 8113 42103 8171 42109
rect 7852 42004 7880 42103
rect 8478 42100 8484 42112
rect 8536 42100 8542 42152
rect 12253 42143 12311 42149
rect 12253 42109 12265 42143
rect 12299 42109 12311 42143
rect 12253 42103 12311 42109
rect 11146 42032 11152 42084
rect 11204 42072 11210 42084
rect 12268 42072 12296 42103
rect 13354 42100 13360 42152
rect 13412 42140 13418 42152
rect 13633 42143 13691 42149
rect 13633 42140 13645 42143
rect 13412 42112 13645 42140
rect 13412 42100 13418 42112
rect 13633 42109 13645 42112
rect 13679 42109 13691 42143
rect 13633 42103 13691 42109
rect 13909 42143 13967 42149
rect 13909 42109 13921 42143
rect 13955 42140 13967 42143
rect 16022 42140 16028 42152
rect 13955 42112 16028 42140
rect 13955 42109 13967 42112
rect 13909 42103 13967 42109
rect 16022 42100 16028 42112
rect 16080 42100 16086 42152
rect 18141 42143 18199 42149
rect 18141 42109 18153 42143
rect 18187 42140 18199 42143
rect 18598 42140 18604 42152
rect 18187 42112 18604 42140
rect 18187 42109 18199 42112
rect 18141 42103 18199 42109
rect 18598 42100 18604 42112
rect 18656 42140 18662 42152
rect 19334 42140 19340 42152
rect 18656 42112 19340 42140
rect 18656 42100 18662 42112
rect 19334 42100 19340 42112
rect 19392 42100 19398 42152
rect 21266 42100 21272 42152
rect 21324 42140 21330 42152
rect 21910 42140 21916 42152
rect 21324 42112 21916 42140
rect 21324 42100 21330 42112
rect 21910 42100 21916 42112
rect 21968 42140 21974 42152
rect 21968 42112 22094 42140
rect 21968 42100 21974 42112
rect 11204 42044 12296 42072
rect 22066 42072 22094 42112
rect 22186 42100 22192 42152
rect 22244 42140 22250 42152
rect 22557 42143 22615 42149
rect 22557 42140 22569 42143
rect 22244 42112 22569 42140
rect 22244 42100 22250 42112
rect 22557 42109 22569 42112
rect 22603 42109 22615 42143
rect 22557 42103 22615 42109
rect 22066 42044 22508 42072
rect 11204 42032 11210 42044
rect 9398 42004 9404 42016
rect 7852 41976 9404 42004
rect 9398 41964 9404 41976
rect 9456 41964 9462 42016
rect 9585 42007 9643 42013
rect 9585 41973 9597 42007
rect 9631 42004 9643 42007
rect 11422 42004 11428 42016
rect 9631 41976 11428 42004
rect 9631 41973 9643 41976
rect 9585 41967 9643 41973
rect 11422 41964 11428 41976
rect 11480 41964 11486 42016
rect 13906 41964 13912 42016
rect 13964 42004 13970 42016
rect 14918 42004 14924 42016
rect 13964 41976 14924 42004
rect 13964 41964 13970 41976
rect 14918 41964 14924 41976
rect 14976 42004 14982 42016
rect 15381 42007 15439 42013
rect 15381 42004 15393 42007
rect 14976 41976 15393 42004
rect 14976 41964 14982 41976
rect 15381 41973 15393 41976
rect 15427 41973 15439 42007
rect 15381 41967 15439 41973
rect 21910 41964 21916 42016
rect 21968 42004 21974 42016
rect 22005 42007 22063 42013
rect 22005 42004 22017 42007
rect 21968 41976 22017 42004
rect 21968 41964 21974 41976
rect 22005 41973 22017 41976
rect 22051 41973 22063 42007
rect 22480 42004 22508 42044
rect 25041 42007 25099 42013
rect 25041 42004 25053 42007
rect 22480 41976 25053 42004
rect 22005 41967 22063 41973
rect 25041 41973 25053 41976
rect 25087 41973 25099 42007
rect 25041 41967 25099 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 3418 41760 3424 41812
rect 3476 41800 3482 41812
rect 4525 41803 4583 41809
rect 4525 41800 4537 41803
rect 3476 41772 4537 41800
rect 3476 41760 3482 41772
rect 4525 41769 4537 41772
rect 4571 41769 4583 41803
rect 4525 41763 4583 41769
rect 7834 41760 7840 41812
rect 7892 41760 7898 41812
rect 17218 41760 17224 41812
rect 17276 41800 17282 41812
rect 25133 41803 25191 41809
rect 25133 41800 25145 41803
rect 17276 41772 25145 41800
rect 17276 41760 17282 41772
rect 25133 41769 25145 41772
rect 25179 41769 25191 41803
rect 25133 41763 25191 41769
rect 5537 41735 5595 41741
rect 5537 41701 5549 41735
rect 5583 41732 5595 41735
rect 5626 41732 5632 41744
rect 5583 41704 5632 41732
rect 5583 41701 5595 41704
rect 5537 41695 5595 41701
rect 5626 41692 5632 41704
rect 5684 41692 5690 41744
rect 19058 41692 19064 41744
rect 19116 41732 19122 41744
rect 19116 41704 20116 41732
rect 19116 41692 19122 41704
rect 8478 41624 8484 41676
rect 8536 41624 8542 41676
rect 11333 41667 11391 41673
rect 11333 41633 11345 41667
rect 11379 41664 11391 41667
rect 11698 41664 11704 41676
rect 11379 41636 11704 41664
rect 11379 41633 11391 41636
rect 11333 41627 11391 41633
rect 11698 41624 11704 41636
rect 11756 41624 11762 41676
rect 13354 41624 13360 41676
rect 13412 41664 13418 41676
rect 15286 41664 15292 41676
rect 13412 41636 15292 41664
rect 13412 41624 13418 41636
rect 15286 41624 15292 41636
rect 15344 41624 15350 41676
rect 17862 41624 17868 41676
rect 17920 41664 17926 41676
rect 18693 41667 18751 41673
rect 18693 41664 18705 41667
rect 17920 41636 18705 41664
rect 17920 41624 17926 41636
rect 18693 41633 18705 41636
rect 18739 41664 18751 41667
rect 18782 41664 18788 41676
rect 18739 41636 18788 41664
rect 18739 41633 18751 41636
rect 18693 41627 18751 41633
rect 18782 41624 18788 41636
rect 18840 41624 18846 41676
rect 19702 41624 19708 41676
rect 19760 41664 19766 41676
rect 20088 41673 20116 41704
rect 20254 41692 20260 41744
rect 20312 41732 20318 41744
rect 24946 41732 24952 41744
rect 20312 41704 24952 41732
rect 20312 41692 20318 41704
rect 24946 41692 24952 41704
rect 25004 41692 25010 41744
rect 19889 41667 19947 41673
rect 19889 41664 19901 41667
rect 19760 41636 19901 41664
rect 19760 41624 19766 41636
rect 19889 41633 19901 41636
rect 19935 41633 19947 41667
rect 19889 41627 19947 41633
rect 20073 41667 20131 41673
rect 20073 41633 20085 41667
rect 20119 41664 20131 41667
rect 21174 41664 21180 41676
rect 20119 41636 21180 41664
rect 20119 41633 20131 41636
rect 20073 41627 20131 41633
rect 21174 41624 21180 41636
rect 21232 41624 21238 41676
rect 21726 41624 21732 41676
rect 21784 41664 21790 41676
rect 22097 41667 22155 41673
rect 22097 41664 22109 41667
rect 21784 41636 22109 41664
rect 21784 41624 21790 41636
rect 22097 41633 22109 41636
rect 22143 41633 22155 41667
rect 22097 41627 22155 41633
rect 4433 41599 4491 41605
rect 4433 41565 4445 41599
rect 4479 41596 4491 41599
rect 6270 41596 6276 41608
rect 4479 41568 6276 41596
rect 4479 41565 4491 41568
rect 4433 41559 4491 41565
rect 6270 41556 6276 41568
rect 6328 41556 6334 41608
rect 8294 41556 8300 41608
rect 8352 41596 8358 41608
rect 10594 41596 10600 41608
rect 8352 41568 10600 41596
rect 8352 41556 8358 41568
rect 10594 41556 10600 41568
rect 10652 41556 10658 41608
rect 17957 41599 18015 41605
rect 17957 41565 17969 41599
rect 18003 41596 18015 41599
rect 19426 41596 19432 41608
rect 18003 41568 19432 41596
rect 18003 41565 18015 41568
rect 17957 41559 18015 41565
rect 19426 41556 19432 41568
rect 19484 41556 19490 41608
rect 21082 41556 21088 41608
rect 21140 41596 21146 41608
rect 21818 41596 21824 41608
rect 21140 41568 21824 41596
rect 21140 41556 21146 41568
rect 21818 41556 21824 41568
rect 21876 41596 21882 41608
rect 21913 41599 21971 41605
rect 21913 41596 21925 41599
rect 21876 41568 21925 41596
rect 21876 41556 21882 41568
rect 21913 41565 21925 41568
rect 21959 41565 21971 41599
rect 21913 41559 21971 41565
rect 22005 41599 22063 41605
rect 22005 41565 22017 41599
rect 22051 41596 22063 41599
rect 22738 41596 22744 41608
rect 22051 41568 22744 41596
rect 22051 41565 22063 41568
rect 22005 41559 22063 41565
rect 22738 41556 22744 41568
rect 22796 41556 22802 41608
rect 23198 41556 23204 41608
rect 23256 41556 23262 41608
rect 23477 41599 23535 41605
rect 23477 41565 23489 41599
rect 23523 41596 23535 41599
rect 23934 41596 23940 41608
rect 23523 41568 23940 41596
rect 23523 41565 23535 41568
rect 23477 41559 23535 41565
rect 23934 41556 23940 41568
rect 23992 41556 23998 41608
rect 25314 41556 25320 41608
rect 25372 41556 25378 41608
rect 1670 41488 1676 41540
rect 1728 41488 1734 41540
rect 1857 41531 1915 41537
rect 1857 41497 1869 41531
rect 1903 41528 1915 41531
rect 3970 41528 3976 41540
rect 1903 41500 3976 41528
rect 1903 41497 1915 41500
rect 1857 41491 1915 41497
rect 3970 41488 3976 41500
rect 4028 41488 4034 41540
rect 5350 41488 5356 41540
rect 5408 41488 5414 41540
rect 11609 41531 11667 41537
rect 11609 41528 11621 41531
rect 11440 41500 11621 41528
rect 11440 41472 11468 41500
rect 11609 41497 11621 41500
rect 11655 41497 11667 41531
rect 11609 41491 11667 41497
rect 12066 41488 12072 41540
rect 12124 41488 12130 41540
rect 15565 41531 15623 41537
rect 15565 41528 15577 41531
rect 13096 41500 15577 41528
rect 7834 41420 7840 41472
rect 7892 41460 7898 41472
rect 8205 41463 8263 41469
rect 8205 41460 8217 41463
rect 7892 41432 8217 41460
rect 7892 41420 7898 41432
rect 8205 41429 8217 41432
rect 8251 41429 8263 41463
rect 8205 41423 8263 41429
rect 8297 41463 8355 41469
rect 8297 41429 8309 41463
rect 8343 41460 8355 41463
rect 9582 41460 9588 41472
rect 8343 41432 9588 41460
rect 8343 41429 8355 41432
rect 8297 41423 8355 41429
rect 9582 41420 9588 41432
rect 9640 41420 9646 41472
rect 11422 41420 11428 41472
rect 11480 41420 11486 41472
rect 12618 41420 12624 41472
rect 12676 41460 12682 41472
rect 13096 41469 13124 41500
rect 15565 41497 15577 41500
rect 15611 41497 15623 41531
rect 18506 41528 18512 41540
rect 15565 41491 15623 41497
rect 15948 41500 16054 41528
rect 16960 41500 18512 41528
rect 13081 41463 13139 41469
rect 13081 41460 13093 41463
rect 12676 41432 13093 41460
rect 12676 41420 12682 41432
rect 13081 41429 13093 41432
rect 13127 41429 13139 41463
rect 13081 41423 13139 41429
rect 14366 41420 14372 41472
rect 14424 41460 14430 41472
rect 15948 41460 15976 41500
rect 16574 41460 16580 41472
rect 14424 41432 16580 41460
rect 14424 41420 14430 41432
rect 16574 41420 16580 41432
rect 16632 41460 16638 41472
rect 16960 41460 16988 41500
rect 18506 41488 18512 41500
rect 18564 41488 18570 41540
rect 16632 41432 16988 41460
rect 17037 41463 17095 41469
rect 16632 41420 16638 41432
rect 17037 41429 17049 41463
rect 17083 41460 17095 41463
rect 18322 41460 18328 41472
rect 17083 41432 18328 41460
rect 17083 41429 17095 41432
rect 17037 41423 17095 41429
rect 18322 41420 18328 41432
rect 18380 41420 18386 41472
rect 19334 41420 19340 41472
rect 19392 41460 19398 41472
rect 19429 41463 19487 41469
rect 19429 41460 19441 41463
rect 19392 41432 19441 41460
rect 19392 41420 19398 41432
rect 19429 41429 19441 41432
rect 19475 41429 19487 41463
rect 19429 41423 19487 41429
rect 19518 41420 19524 41472
rect 19576 41460 19582 41472
rect 19797 41463 19855 41469
rect 19797 41460 19809 41463
rect 19576 41432 19809 41460
rect 19576 41420 19582 41432
rect 19797 41429 19809 41432
rect 19843 41429 19855 41463
rect 19797 41423 19855 41429
rect 21542 41420 21548 41472
rect 21600 41420 21606 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 3510 41216 3516 41268
rect 3568 41256 3574 41268
rect 4065 41259 4123 41265
rect 4065 41256 4077 41259
rect 3568 41228 4077 41256
rect 3568 41216 3574 41228
rect 4065 41225 4077 41228
rect 4111 41225 4123 41259
rect 4065 41219 4123 41225
rect 7006 41216 7012 41268
rect 7064 41256 7070 41268
rect 7558 41256 7564 41268
rect 7064 41228 7564 41256
rect 7064 41216 7070 41228
rect 7558 41216 7564 41228
rect 7616 41216 7622 41268
rect 8297 41259 8355 41265
rect 8297 41225 8309 41259
rect 8343 41256 8355 41259
rect 8478 41256 8484 41268
rect 8343 41228 8484 41256
rect 8343 41225 8355 41228
rect 8297 41219 8355 41225
rect 8478 41216 8484 41228
rect 8536 41216 8542 41268
rect 11701 41259 11759 41265
rect 10060 41228 11652 41256
rect 10060 41188 10088 41228
rect 11624 41188 11652 41228
rect 11701 41225 11713 41259
rect 11747 41256 11759 41259
rect 11974 41256 11980 41268
rect 11747 41228 11980 41256
rect 11747 41225 11759 41228
rect 11701 41219 11759 41225
rect 11974 41216 11980 41228
rect 12032 41216 12038 41268
rect 12066 41216 12072 41268
rect 12124 41216 12130 41268
rect 12161 41259 12219 41265
rect 12161 41225 12173 41259
rect 12207 41256 12219 41259
rect 15102 41256 15108 41268
rect 12207 41228 15108 41256
rect 12207 41225 12219 41228
rect 12161 41219 12219 41225
rect 15102 41216 15108 41228
rect 15160 41216 15166 41268
rect 17310 41216 17316 41268
rect 17368 41216 17374 41268
rect 20806 41256 20812 41268
rect 18340 41228 20812 41256
rect 12084 41188 12112 41216
rect 8312 41160 10166 41188
rect 11624 41160 12112 41188
rect 13633 41191 13691 41197
rect 8312 41132 8340 41160
rect 13633 41157 13645 41191
rect 13679 41188 13691 41191
rect 13906 41188 13912 41200
rect 13679 41160 13912 41188
rect 13679 41157 13691 41160
rect 13633 41151 13691 41157
rect 13906 41148 13912 41160
rect 13964 41148 13970 41200
rect 14274 41148 14280 41200
rect 14332 41148 14338 41200
rect 17221 41191 17279 41197
rect 17221 41157 17233 41191
rect 17267 41188 17279 41191
rect 18340 41188 18368 41228
rect 20806 41216 20812 41228
rect 20864 41256 20870 41268
rect 21450 41256 21456 41268
rect 20864 41228 21456 41256
rect 20864 41216 20870 41228
rect 21450 41216 21456 41228
rect 21508 41216 21514 41268
rect 22465 41259 22523 41265
rect 22465 41225 22477 41259
rect 22511 41256 22523 41259
rect 22830 41256 22836 41268
rect 22511 41228 22836 41256
rect 22511 41225 22523 41228
rect 22465 41219 22523 41225
rect 22830 41216 22836 41228
rect 22888 41216 22894 41268
rect 18782 41188 18788 41200
rect 17267 41160 18368 41188
rect 18432 41160 18788 41188
rect 17267 41157 17279 41160
rect 17221 41151 17279 41157
rect 3973 41123 4031 41129
rect 3973 41089 3985 41123
rect 4019 41120 4031 41123
rect 4062 41120 4068 41132
rect 4019 41092 4068 41120
rect 4019 41089 4031 41092
rect 3973 41083 4031 41089
rect 4062 41080 4068 41092
rect 4120 41080 4126 41132
rect 8294 41120 8300 41132
rect 7958 41092 8300 41120
rect 8294 41080 8300 41092
rect 8352 41080 8358 41132
rect 12066 41080 12072 41132
rect 12124 41080 12130 41132
rect 13354 41080 13360 41132
rect 13412 41080 13418 41132
rect 18432 41129 18460 41160
rect 18782 41148 18788 41160
rect 18840 41148 18846 41200
rect 19242 41148 19248 41200
rect 19300 41148 19306 41200
rect 21082 41148 21088 41200
rect 21140 41188 21146 41200
rect 22002 41188 22008 41200
rect 21140 41160 22008 41188
rect 21140 41148 21146 41160
rect 22002 41148 22008 41160
rect 22060 41188 22066 41200
rect 22060 41160 23244 41188
rect 22060 41148 22066 41160
rect 18417 41123 18475 41129
rect 18417 41089 18429 41123
rect 18463 41089 18475 41123
rect 18417 41083 18475 41089
rect 22094 41080 22100 41132
rect 22152 41120 22158 41132
rect 23216 41129 23244 41160
rect 23474 41148 23480 41200
rect 23532 41148 23538 41200
rect 24486 41148 24492 41200
rect 24544 41148 24550 41200
rect 22373 41123 22431 41129
rect 22373 41120 22385 41123
rect 22152 41092 22385 41120
rect 22152 41080 22158 41092
rect 22373 41089 22385 41092
rect 22419 41089 22431 41123
rect 22373 41083 22431 41089
rect 23201 41123 23259 41129
rect 23201 41089 23213 41123
rect 23247 41089 23259 41123
rect 23201 41083 23259 41089
rect 6270 41012 6276 41064
rect 6328 41052 6334 41064
rect 6549 41055 6607 41061
rect 6549 41052 6561 41055
rect 6328 41024 6561 41052
rect 6328 41012 6334 41024
rect 6549 41021 6561 41024
rect 6595 41021 6607 41055
rect 6549 41015 6607 41021
rect 6825 41055 6883 41061
rect 6825 41021 6837 41055
rect 6871 41052 6883 41055
rect 7558 41052 7564 41064
rect 6871 41024 7564 41052
rect 6871 41021 6883 41024
rect 6825 41015 6883 41021
rect 6564 40916 6592 41015
rect 7558 41012 7564 41024
rect 7616 41012 7622 41064
rect 9398 41052 9404 41064
rect 7852 41024 9404 41052
rect 7852 40916 7880 41024
rect 9398 41012 9404 41024
rect 9456 41012 9462 41064
rect 9677 41055 9735 41061
rect 9677 41021 9689 41055
rect 9723 41052 9735 41055
rect 11606 41052 11612 41064
rect 9723 41024 11612 41052
rect 9723 41021 9735 41024
rect 9677 41015 9735 41021
rect 11606 41012 11612 41024
rect 11664 41012 11670 41064
rect 12342 41012 12348 41064
rect 12400 41012 12406 41064
rect 13998 41012 14004 41064
rect 14056 41052 14062 41064
rect 17405 41055 17463 41061
rect 17405 41052 17417 41055
rect 14056 41024 17417 41052
rect 14056 41012 14062 41024
rect 17405 41021 17417 41024
rect 17451 41021 17463 41055
rect 17405 41015 17463 41021
rect 18690 41012 18696 41064
rect 18748 41052 18754 41064
rect 19058 41052 19064 41064
rect 18748 41024 19064 41052
rect 18748 41012 18754 41024
rect 19058 41012 19064 41024
rect 19116 41012 19122 41064
rect 22554 41012 22560 41064
rect 22612 41052 22618 41064
rect 22649 41055 22707 41061
rect 22649 41052 22661 41055
rect 22612 41024 22661 41052
rect 22612 41012 22618 41024
rect 22649 41021 22661 41024
rect 22695 41052 22707 41055
rect 22695 41024 24992 41052
rect 22695 41021 22707 41024
rect 22649 41015 22707 41021
rect 6564 40888 7880 40916
rect 11146 40876 11152 40928
rect 11204 40876 11210 40928
rect 14918 40876 14924 40928
rect 14976 40916 14982 40928
rect 15105 40919 15163 40925
rect 15105 40916 15117 40919
rect 14976 40888 15117 40916
rect 14976 40876 14982 40888
rect 15105 40885 15117 40888
rect 15151 40885 15163 40919
rect 15105 40879 15163 40885
rect 16850 40876 16856 40928
rect 16908 40876 16914 40928
rect 18506 40876 18512 40928
rect 18564 40916 18570 40928
rect 18782 40916 18788 40928
rect 18564 40888 18788 40916
rect 18564 40876 18570 40888
rect 18782 40876 18788 40888
rect 18840 40916 18846 40928
rect 19242 40916 19248 40928
rect 18840 40888 19248 40916
rect 18840 40876 18846 40888
rect 19242 40876 19248 40888
rect 19300 40876 19306 40928
rect 20070 40876 20076 40928
rect 20128 40916 20134 40928
rect 20165 40919 20223 40925
rect 20165 40916 20177 40919
rect 20128 40888 20177 40916
rect 20128 40876 20134 40888
rect 20165 40885 20177 40888
rect 20211 40885 20223 40919
rect 20165 40879 20223 40885
rect 21450 40876 21456 40928
rect 21508 40876 21514 40928
rect 22005 40919 22063 40925
rect 22005 40885 22017 40919
rect 22051 40916 22063 40919
rect 23658 40916 23664 40928
rect 22051 40888 23664 40916
rect 22051 40885 22063 40888
rect 22005 40879 22063 40885
rect 23658 40876 23664 40888
rect 23716 40876 23722 40928
rect 24964 40925 24992 41024
rect 24949 40919 25007 40925
rect 24949 40885 24961 40919
rect 24995 40916 25007 40919
rect 25038 40916 25044 40928
rect 24995 40888 25044 40916
rect 24995 40885 25007 40888
rect 24949 40879 25007 40885
rect 25038 40876 25044 40888
rect 25096 40876 25102 40928
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 1578 40672 1584 40724
rect 1636 40712 1642 40724
rect 2869 40715 2927 40721
rect 2869 40712 2881 40715
rect 1636 40684 2881 40712
rect 1636 40672 1642 40684
rect 2869 40681 2881 40684
rect 2915 40681 2927 40715
rect 2869 40675 2927 40681
rect 15194 40672 15200 40724
rect 15252 40712 15258 40724
rect 17313 40715 17371 40721
rect 17313 40712 17325 40715
rect 15252 40684 17325 40712
rect 15252 40672 15258 40684
rect 17313 40681 17325 40684
rect 17359 40681 17371 40715
rect 17313 40675 17371 40681
rect 17678 40672 17684 40724
rect 17736 40712 17742 40724
rect 17862 40712 17868 40724
rect 17736 40684 17868 40712
rect 17736 40672 17742 40684
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 21358 40712 21364 40724
rect 21008 40684 21364 40712
rect 12805 40647 12863 40653
rect 12805 40613 12817 40647
rect 12851 40644 12863 40647
rect 13814 40644 13820 40656
rect 12851 40616 13820 40644
rect 12851 40613 12863 40616
rect 12805 40607 12863 40613
rect 13814 40604 13820 40616
rect 13872 40604 13878 40656
rect 15841 40647 15899 40653
rect 15841 40613 15853 40647
rect 15887 40644 15899 40647
rect 19058 40644 19064 40656
rect 15887 40616 19064 40644
rect 15887 40613 15899 40616
rect 15841 40607 15899 40613
rect 19058 40604 19064 40616
rect 19116 40604 19122 40656
rect 12158 40536 12164 40588
rect 12216 40576 12222 40588
rect 12216 40548 12434 40576
rect 12216 40536 12222 40548
rect 6270 40468 6276 40520
rect 6328 40468 6334 40520
rect 12406 40452 12434 40548
rect 12618 40536 12624 40588
rect 12676 40576 12682 40588
rect 13357 40579 13415 40585
rect 13357 40576 13369 40579
rect 12676 40548 13369 40576
rect 12676 40536 12682 40548
rect 13357 40545 13369 40548
rect 13403 40545 13415 40579
rect 13357 40539 13415 40545
rect 16390 40536 16396 40588
rect 16448 40536 16454 40588
rect 16482 40536 16488 40588
rect 16540 40576 16546 40588
rect 17865 40579 17923 40585
rect 17865 40576 17877 40579
rect 16540 40548 17877 40576
rect 16540 40536 16546 40548
rect 17865 40545 17877 40548
rect 17911 40545 17923 40579
rect 17865 40539 17923 40545
rect 18598 40536 18604 40588
rect 18656 40536 18662 40588
rect 19610 40536 19616 40588
rect 19668 40576 19674 40588
rect 19889 40579 19947 40585
rect 19889 40576 19901 40579
rect 19668 40548 19901 40576
rect 19668 40536 19674 40548
rect 19889 40545 19901 40548
rect 19935 40545 19947 40579
rect 19889 40539 19947 40545
rect 19981 40579 20039 40585
rect 19981 40545 19993 40579
rect 20027 40545 20039 40579
rect 19981 40539 20039 40545
rect 13173 40511 13231 40517
rect 13173 40477 13185 40511
rect 13219 40508 13231 40511
rect 13446 40508 13452 40520
rect 13219 40480 13452 40508
rect 13219 40477 13231 40480
rect 13173 40471 13231 40477
rect 13446 40468 13452 40480
rect 13504 40468 13510 40520
rect 16301 40511 16359 40517
rect 16301 40477 16313 40511
rect 16347 40508 16359 40511
rect 16666 40508 16672 40520
rect 16347 40480 16672 40508
rect 16347 40477 16359 40480
rect 16301 40471 16359 40477
rect 16666 40468 16672 40480
rect 16724 40468 16730 40520
rect 18322 40468 18328 40520
rect 18380 40468 18386 40520
rect 18506 40468 18512 40520
rect 18564 40508 18570 40520
rect 18616 40508 18644 40536
rect 19996 40508 20024 40539
rect 18564 40480 20024 40508
rect 18564 40468 18570 40480
rect 2777 40443 2835 40449
rect 2777 40409 2789 40443
rect 2823 40440 2835 40443
rect 5074 40440 5080 40452
rect 2823 40412 5080 40440
rect 2823 40409 2835 40412
rect 2777 40403 2835 40409
rect 5074 40400 5080 40412
rect 5132 40400 5138 40452
rect 6546 40400 6552 40452
rect 6604 40400 6610 40452
rect 8294 40440 8300 40452
rect 7774 40412 8300 40440
rect 8294 40400 8300 40412
rect 8352 40400 8358 40452
rect 11422 40400 11428 40452
rect 11480 40400 11486 40452
rect 11790 40400 11796 40452
rect 11848 40440 11854 40452
rect 12158 40440 12164 40452
rect 11848 40412 12164 40440
rect 11848 40400 11854 40412
rect 12158 40400 12164 40412
rect 12216 40400 12222 40452
rect 12342 40400 12348 40452
rect 12400 40440 12434 40452
rect 14274 40440 14280 40452
rect 12400 40412 14280 40440
rect 12400 40400 12406 40412
rect 14274 40400 14280 40412
rect 14332 40400 14338 40452
rect 18340 40440 18368 40468
rect 18598 40440 18604 40452
rect 18340 40412 18604 40440
rect 18598 40400 18604 40412
rect 18656 40400 18662 40452
rect 19797 40443 19855 40449
rect 19797 40409 19809 40443
rect 19843 40440 19855 40443
rect 21008 40440 21036 40684
rect 21358 40672 21364 40684
rect 21416 40672 21422 40724
rect 21082 40536 21088 40588
rect 21140 40536 21146 40588
rect 23566 40536 23572 40588
rect 23624 40576 23630 40588
rect 23845 40579 23903 40585
rect 23845 40576 23857 40579
rect 23624 40548 23857 40576
rect 23624 40536 23630 40548
rect 23845 40545 23857 40548
rect 23891 40545 23903 40579
rect 23845 40539 23903 40545
rect 23658 40468 23664 40520
rect 23716 40508 23722 40520
rect 23753 40511 23811 40517
rect 23753 40508 23765 40511
rect 23716 40480 23765 40508
rect 23716 40468 23722 40480
rect 23753 40477 23765 40480
rect 23799 40477 23811 40511
rect 23753 40471 23811 40477
rect 24765 40511 24823 40517
rect 24765 40477 24777 40511
rect 24811 40508 24823 40511
rect 24946 40508 24952 40520
rect 24811 40480 24952 40508
rect 24811 40477 24823 40480
rect 24765 40471 24823 40477
rect 24946 40468 24952 40480
rect 25004 40468 25010 40520
rect 19843 40412 21036 40440
rect 19843 40409 19855 40412
rect 19797 40403 19855 40409
rect 21266 40400 21272 40452
rect 21324 40440 21330 40452
rect 21361 40443 21419 40449
rect 21361 40440 21373 40443
rect 21324 40412 21373 40440
rect 21324 40400 21330 40412
rect 21361 40409 21373 40412
rect 21407 40409 21419 40443
rect 24394 40440 24400 40452
rect 22586 40412 24400 40440
rect 21361 40403 21419 40409
rect 24394 40400 24400 40412
rect 24452 40400 24458 40452
rect 7558 40332 7564 40384
rect 7616 40372 7622 40384
rect 8021 40375 8079 40381
rect 8021 40372 8033 40375
rect 7616 40344 8033 40372
rect 7616 40332 7622 40344
rect 8021 40341 8033 40344
rect 8067 40341 8079 40375
rect 8021 40335 8079 40341
rect 13265 40375 13323 40381
rect 13265 40341 13277 40375
rect 13311 40372 13323 40375
rect 15746 40372 15752 40384
rect 13311 40344 15752 40372
rect 13311 40341 13323 40344
rect 13265 40335 13323 40341
rect 15746 40332 15752 40344
rect 15804 40332 15810 40384
rect 16206 40332 16212 40384
rect 16264 40332 16270 40384
rect 17678 40332 17684 40384
rect 17736 40332 17742 40384
rect 17773 40375 17831 40381
rect 17773 40341 17785 40375
rect 17819 40372 17831 40375
rect 18322 40372 18328 40384
rect 17819 40344 18328 40372
rect 17819 40341 17831 40344
rect 17773 40335 17831 40341
rect 18322 40332 18328 40344
rect 18380 40332 18386 40384
rect 19429 40375 19487 40381
rect 19429 40341 19441 40375
rect 19475 40372 19487 40375
rect 19702 40372 19708 40384
rect 19475 40344 19708 40372
rect 19475 40341 19487 40344
rect 19429 40335 19487 40341
rect 19702 40332 19708 40344
rect 19760 40332 19766 40384
rect 22830 40332 22836 40384
rect 22888 40332 22894 40384
rect 23293 40375 23351 40381
rect 23293 40341 23305 40375
rect 23339 40372 23351 40375
rect 23566 40372 23572 40384
rect 23339 40344 23572 40372
rect 23339 40341 23351 40344
rect 23293 40335 23351 40341
rect 23566 40332 23572 40344
rect 23624 40332 23630 40384
rect 23658 40332 23664 40384
rect 23716 40332 23722 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7837 40171 7895 40177
rect 7837 40137 7849 40171
rect 7883 40168 7895 40171
rect 8754 40168 8760 40180
rect 7883 40140 8760 40168
rect 7883 40137 7895 40140
rect 7837 40131 7895 40137
rect 8754 40128 8760 40140
rect 8812 40128 8818 40180
rect 11422 40168 11428 40180
rect 9048 40140 11428 40168
rect 6086 40060 6092 40112
rect 6144 40100 6150 40112
rect 9048 40109 9076 40140
rect 11422 40128 11428 40140
rect 11480 40128 11486 40180
rect 12526 40168 12532 40180
rect 12176 40140 12532 40168
rect 8205 40103 8263 40109
rect 8205 40100 8217 40103
rect 6144 40072 8217 40100
rect 6144 40060 6150 40072
rect 8205 40069 8217 40072
rect 8251 40100 8263 40103
rect 9033 40103 9091 40109
rect 8251 40072 8984 40100
rect 8251 40069 8263 40072
rect 8205 40063 8263 40069
rect 3878 39992 3884 40044
rect 3936 40032 3942 40044
rect 8297 40035 8355 40041
rect 8297 40032 8309 40035
rect 3936 40004 8309 40032
rect 3936 39992 3942 40004
rect 8297 40001 8309 40004
rect 8343 40032 8355 40035
rect 8956 40032 8984 40072
rect 9033 40069 9045 40103
rect 9079 40069 9091 40103
rect 9033 40063 9091 40069
rect 9398 40060 9404 40112
rect 9456 40100 9462 40112
rect 9769 40103 9827 40109
rect 9769 40100 9781 40103
rect 9456 40072 9781 40100
rect 9456 40060 9462 40072
rect 9769 40069 9781 40072
rect 9815 40069 9827 40103
rect 9769 40063 9827 40069
rect 9858 40032 9864 40044
rect 8343 40004 8892 40032
rect 8956 40004 9864 40032
rect 8343 40001 8355 40004
rect 8297 39995 8355 40001
rect 8389 39967 8447 39973
rect 8389 39933 8401 39967
rect 8435 39933 8447 39967
rect 8864 39964 8892 40004
rect 9858 39992 9864 40004
rect 9916 39992 9922 40044
rect 12176 40032 12204 40140
rect 12526 40128 12532 40140
rect 12584 40128 12590 40180
rect 20717 40171 20775 40177
rect 20717 40137 20729 40171
rect 20763 40137 20775 40171
rect 20717 40131 20775 40137
rect 21085 40171 21143 40177
rect 21085 40137 21097 40171
rect 21131 40168 21143 40171
rect 21450 40168 21456 40180
rect 21131 40140 21456 40168
rect 21131 40137 21143 40140
rect 21085 40131 21143 40137
rect 12434 40060 12440 40112
rect 12492 40100 12498 40112
rect 12492 40072 12926 40100
rect 12492 40060 12498 40072
rect 13906 40060 13912 40112
rect 13964 40100 13970 40112
rect 14274 40100 14280 40112
rect 13964 40072 14280 40100
rect 13964 40060 13970 40072
rect 14274 40060 14280 40072
rect 14332 40060 14338 40112
rect 15565 40103 15623 40109
rect 15565 40069 15577 40103
rect 15611 40100 15623 40103
rect 20254 40100 20260 40112
rect 15611 40072 20260 40100
rect 15611 40069 15623 40072
rect 15565 40063 15623 40069
rect 20254 40060 20260 40072
rect 20312 40060 20318 40112
rect 20732 40100 20760 40131
rect 21450 40128 21456 40140
rect 21508 40128 21514 40180
rect 22005 40171 22063 40177
rect 22005 40137 22017 40171
rect 22051 40168 22063 40171
rect 23842 40168 23848 40180
rect 22051 40140 23848 40168
rect 22051 40137 22063 40140
rect 22005 40131 22063 40137
rect 23842 40128 23848 40140
rect 23900 40128 23906 40180
rect 22373 40103 22431 40109
rect 22373 40100 22385 40103
rect 20732 40072 22385 40100
rect 22373 40069 22385 40072
rect 22419 40069 22431 40103
rect 22373 40063 22431 40069
rect 12084 40004 12204 40032
rect 12084 39964 12112 40004
rect 21910 39992 21916 40044
rect 21968 40032 21974 40044
rect 22465 40035 22523 40041
rect 22465 40032 22477 40035
rect 21968 40004 22477 40032
rect 21968 39992 21974 40004
rect 22465 40001 22477 40004
rect 22511 40001 22523 40035
rect 22465 39995 22523 40001
rect 23201 40035 23259 40041
rect 23201 40001 23213 40035
rect 23247 40032 23259 40035
rect 24854 40032 24860 40044
rect 23247 40004 24860 40032
rect 23247 40001 23259 40004
rect 23201 39995 23259 40001
rect 24854 39992 24860 40004
rect 24912 39992 24918 40044
rect 8864 39936 12112 39964
rect 8389 39927 8447 39933
rect 7282 39856 7288 39908
rect 7340 39896 7346 39908
rect 8404 39896 8432 39927
rect 12158 39924 12164 39976
rect 12216 39924 12222 39976
rect 12434 39924 12440 39976
rect 12492 39924 12498 39976
rect 12526 39924 12532 39976
rect 12584 39964 12590 39976
rect 15010 39964 15016 39976
rect 12584 39936 15016 39964
rect 12584 39924 12590 39936
rect 15010 39924 15016 39936
rect 15068 39964 15074 39976
rect 15657 39967 15715 39973
rect 15657 39964 15669 39967
rect 15068 39936 15669 39964
rect 15068 39924 15074 39936
rect 15657 39933 15669 39936
rect 15703 39933 15715 39967
rect 15657 39927 15715 39933
rect 15749 39967 15807 39973
rect 15749 39933 15761 39967
rect 15795 39933 15807 39967
rect 15749 39927 15807 39933
rect 7340 39868 8432 39896
rect 7340 39856 7346 39868
rect 9858 39856 9864 39908
rect 9916 39896 9922 39908
rect 11698 39896 11704 39908
rect 9916 39868 11704 39896
rect 9916 39856 9922 39868
rect 11698 39856 11704 39868
rect 11756 39856 11762 39908
rect 13538 39856 13544 39908
rect 13596 39896 13602 39908
rect 15764 39896 15792 39927
rect 17862 39924 17868 39976
rect 17920 39964 17926 39976
rect 19610 39964 19616 39976
rect 17920 39936 19616 39964
rect 17920 39924 17926 39936
rect 19610 39924 19616 39936
rect 19668 39924 19674 39976
rect 21174 39924 21180 39976
rect 21232 39924 21238 39976
rect 21361 39967 21419 39973
rect 21361 39933 21373 39967
rect 21407 39964 21419 39967
rect 22186 39964 22192 39976
rect 21407 39936 22192 39964
rect 21407 39933 21419 39936
rect 21361 39927 21419 39933
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 22278 39924 22284 39976
rect 22336 39964 22342 39976
rect 22557 39967 22615 39973
rect 22557 39964 22569 39967
rect 22336 39936 22569 39964
rect 22336 39924 22342 39936
rect 22557 39933 22569 39936
rect 22603 39933 22615 39967
rect 22557 39927 22615 39933
rect 23477 39967 23535 39973
rect 23477 39933 23489 39967
rect 23523 39933 23535 39967
rect 23477 39927 23535 39933
rect 24489 39967 24547 39973
rect 24489 39933 24501 39967
rect 24535 39933 24547 39967
rect 24489 39927 24547 39933
rect 13596 39868 15792 39896
rect 13596 39856 13602 39868
rect 16574 39856 16580 39908
rect 16632 39896 16638 39908
rect 16632 39868 18920 39896
rect 16632 39856 16638 39868
rect 6546 39788 6552 39840
rect 6604 39828 6610 39840
rect 11238 39828 11244 39840
rect 6604 39800 11244 39828
rect 6604 39788 6610 39800
rect 11238 39788 11244 39800
rect 11296 39788 11302 39840
rect 11606 39788 11612 39840
rect 11664 39828 11670 39840
rect 13906 39828 13912 39840
rect 11664 39800 13912 39828
rect 11664 39788 11670 39800
rect 13906 39788 13912 39800
rect 13964 39788 13970 39840
rect 13998 39788 14004 39840
rect 14056 39828 14062 39840
rect 14553 39831 14611 39837
rect 14553 39828 14565 39831
rect 14056 39800 14565 39828
rect 14056 39788 14062 39800
rect 14553 39797 14565 39800
rect 14599 39797 14611 39831
rect 14553 39791 14611 39797
rect 15194 39788 15200 39840
rect 15252 39788 15258 39840
rect 17494 39788 17500 39840
rect 17552 39828 17558 39840
rect 18046 39828 18052 39840
rect 17552 39800 18052 39828
rect 17552 39788 17558 39800
rect 18046 39788 18052 39800
rect 18104 39788 18110 39840
rect 18414 39788 18420 39840
rect 18472 39828 18478 39840
rect 18782 39828 18788 39840
rect 18472 39800 18788 39828
rect 18472 39788 18478 39800
rect 18782 39788 18788 39800
rect 18840 39788 18846 39840
rect 18892 39828 18920 39868
rect 20530 39856 20536 39908
rect 20588 39896 20594 39908
rect 23492 39896 23520 39927
rect 20588 39868 23520 39896
rect 24504 39896 24532 39927
rect 25130 39896 25136 39908
rect 24504 39868 25136 39896
rect 20588 39856 20594 39868
rect 25130 39856 25136 39868
rect 25188 39856 25194 39908
rect 24719 39831 24777 39837
rect 24719 39828 24731 39831
rect 18892 39800 24731 39828
rect 24719 39797 24731 39800
rect 24765 39797 24777 39831
rect 24719 39791 24777 39797
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 6914 39584 6920 39636
rect 6972 39624 6978 39636
rect 7190 39624 7196 39636
rect 6972 39596 7196 39624
rect 6972 39584 6978 39596
rect 7190 39584 7196 39596
rect 7248 39584 7254 39636
rect 7650 39584 7656 39636
rect 7708 39584 7714 39636
rect 10584 39627 10642 39633
rect 10584 39593 10596 39627
rect 10630 39624 10642 39627
rect 11146 39624 11152 39636
rect 10630 39596 11152 39624
rect 10630 39593 10642 39596
rect 10584 39587 10642 39593
rect 11146 39584 11152 39596
rect 11204 39584 11210 39636
rect 11238 39584 11244 39636
rect 11296 39624 11302 39636
rect 11296 39596 13216 39624
rect 11296 39584 11302 39596
rect 9125 39559 9183 39565
rect 9125 39525 9137 39559
rect 9171 39556 9183 39559
rect 9858 39556 9864 39568
rect 9171 39528 9864 39556
rect 9171 39525 9183 39528
rect 9125 39519 9183 39525
rect 9858 39516 9864 39528
rect 9916 39516 9922 39568
rect 11698 39516 11704 39568
rect 11756 39556 11762 39568
rect 11756 39528 13124 39556
rect 11756 39516 11762 39528
rect 6914 39448 6920 39500
rect 6972 39488 6978 39500
rect 8205 39491 8263 39497
rect 8205 39488 8217 39491
rect 6972 39460 8217 39488
rect 6972 39448 6978 39460
rect 8205 39457 8217 39460
rect 8251 39457 8263 39491
rect 8205 39451 8263 39457
rect 9030 39448 9036 39500
rect 9088 39488 9094 39500
rect 9677 39491 9735 39497
rect 9677 39488 9689 39491
rect 9088 39460 9689 39488
rect 9088 39448 9094 39460
rect 9677 39457 9689 39460
rect 9723 39457 9735 39491
rect 9677 39451 9735 39457
rect 10321 39491 10379 39497
rect 10321 39457 10333 39491
rect 10367 39488 10379 39491
rect 12158 39488 12164 39500
rect 10367 39460 12164 39488
rect 10367 39457 10379 39460
rect 10321 39451 10379 39457
rect 12158 39448 12164 39460
rect 12216 39448 12222 39500
rect 12434 39448 12440 39500
rect 12492 39488 12498 39500
rect 13096 39497 13124 39528
rect 13188 39497 13216 39596
rect 13630 39584 13636 39636
rect 13688 39624 13694 39636
rect 15749 39627 15807 39633
rect 15749 39624 15761 39627
rect 13688 39596 15761 39624
rect 13688 39584 13694 39596
rect 15749 39593 15761 39596
rect 15795 39593 15807 39627
rect 15749 39587 15807 39593
rect 16390 39584 16396 39636
rect 16448 39624 16454 39636
rect 18782 39624 18788 39636
rect 16448 39596 18788 39624
rect 16448 39584 16454 39596
rect 18782 39584 18788 39596
rect 18840 39584 18846 39636
rect 19518 39584 19524 39636
rect 19576 39584 19582 39636
rect 20714 39584 20720 39636
rect 20772 39584 20778 39636
rect 23658 39584 23664 39636
rect 23716 39624 23722 39636
rect 24581 39627 24639 39633
rect 24581 39624 24593 39627
rect 23716 39596 24593 39624
rect 23716 39584 23722 39596
rect 24581 39593 24593 39596
rect 24627 39593 24639 39627
rect 24581 39587 24639 39593
rect 19242 39556 19248 39568
rect 17236 39528 19248 39556
rect 13081 39491 13139 39497
rect 12492 39460 13032 39488
rect 12492 39448 12498 39460
rect 7466 39380 7472 39432
rect 7524 39420 7530 39432
rect 9490 39420 9496 39432
rect 7524 39392 9496 39420
rect 7524 39380 7530 39392
rect 9490 39380 9496 39392
rect 9548 39380 9554 39432
rect 12342 39420 12348 39432
rect 11730 39392 12348 39420
rect 12342 39380 12348 39392
rect 12400 39380 12406 39432
rect 12526 39380 12532 39432
rect 12584 39420 12590 39432
rect 12710 39420 12716 39432
rect 12584 39392 12716 39420
rect 12584 39380 12590 39392
rect 12710 39380 12716 39392
rect 12768 39380 12774 39432
rect 13004 39420 13032 39460
rect 13081 39457 13093 39491
rect 13127 39457 13139 39491
rect 13081 39451 13139 39457
rect 13173 39491 13231 39497
rect 13173 39457 13185 39491
rect 13219 39457 13231 39491
rect 13173 39451 13231 39457
rect 13906 39448 13912 39500
rect 13964 39488 13970 39500
rect 14829 39491 14887 39497
rect 14829 39488 14841 39491
rect 13964 39460 14841 39488
rect 13964 39448 13970 39460
rect 14829 39457 14841 39460
rect 14875 39457 14887 39491
rect 14829 39451 14887 39457
rect 16390 39448 16396 39500
rect 16448 39448 16454 39500
rect 13538 39420 13544 39432
rect 13004 39392 13544 39420
rect 13538 39380 13544 39392
rect 13596 39380 13602 39432
rect 14737 39423 14795 39429
rect 14737 39389 14749 39423
rect 14783 39420 14795 39423
rect 15194 39420 15200 39432
rect 14783 39392 15200 39420
rect 14783 39389 14795 39392
rect 14737 39383 14795 39389
rect 15194 39380 15200 39392
rect 15252 39380 15258 39432
rect 16209 39423 16267 39429
rect 16209 39389 16221 39423
rect 16255 39420 16267 39423
rect 17236 39420 17264 39528
rect 19242 39516 19248 39528
rect 19300 39516 19306 39568
rect 21818 39516 21824 39568
rect 21876 39556 21882 39568
rect 25774 39556 25780 39568
rect 21876 39528 25780 39556
rect 21876 39516 21882 39528
rect 25774 39516 25780 39528
rect 25832 39516 25838 39568
rect 16255 39392 17264 39420
rect 17328 39460 17540 39488
rect 16255 39389 16267 39392
rect 16209 39383 16267 39389
rect 9585 39355 9643 39361
rect 9585 39321 9597 39355
rect 9631 39352 9643 39355
rect 9674 39352 9680 39364
rect 9631 39324 9680 39352
rect 9631 39321 9643 39324
rect 9585 39315 9643 39321
rect 9674 39312 9680 39324
rect 9732 39312 9738 39364
rect 12250 39312 12256 39364
rect 12308 39352 12314 39364
rect 14645 39355 14703 39361
rect 12308 39324 13676 39352
rect 12308 39312 12314 39324
rect 7650 39244 7656 39296
rect 7708 39284 7714 39296
rect 8021 39287 8079 39293
rect 8021 39284 8033 39287
rect 7708 39256 8033 39284
rect 7708 39244 7714 39256
rect 8021 39253 8033 39256
rect 8067 39253 8079 39287
rect 8021 39247 8079 39253
rect 8113 39287 8171 39293
rect 8113 39253 8125 39287
rect 8159 39284 8171 39287
rect 9398 39284 9404 39296
rect 8159 39256 9404 39284
rect 8159 39253 8171 39256
rect 8113 39247 8171 39253
rect 9398 39244 9404 39256
rect 9456 39244 9462 39296
rect 12069 39287 12127 39293
rect 12069 39253 12081 39287
rect 12115 39284 12127 39287
rect 12158 39284 12164 39296
rect 12115 39256 12164 39284
rect 12115 39253 12127 39256
rect 12069 39247 12127 39253
rect 12158 39244 12164 39256
rect 12216 39244 12222 39296
rect 12342 39244 12348 39296
rect 12400 39284 12406 39296
rect 12621 39287 12679 39293
rect 12621 39284 12633 39287
rect 12400 39256 12633 39284
rect 12400 39244 12406 39256
rect 12621 39253 12633 39256
rect 12667 39253 12679 39287
rect 12621 39247 12679 39253
rect 12986 39244 12992 39296
rect 13044 39244 13050 39296
rect 13648 39284 13676 39324
rect 14645 39321 14657 39355
rect 14691 39352 14703 39355
rect 17328 39352 17356 39460
rect 17402 39380 17408 39432
rect 17460 39380 17466 39432
rect 14691 39324 17356 39352
rect 14691 39321 14703 39324
rect 14645 39315 14703 39321
rect 14277 39287 14335 39293
rect 14277 39284 14289 39287
rect 13648 39256 14289 39284
rect 14277 39253 14289 39256
rect 14323 39253 14335 39287
rect 14277 39247 14335 39253
rect 15562 39244 15568 39296
rect 15620 39284 15626 39296
rect 17420 39293 17448 39380
rect 16117 39287 16175 39293
rect 16117 39284 16129 39287
rect 15620 39256 16129 39284
rect 15620 39244 15626 39256
rect 16117 39253 16129 39256
rect 16163 39253 16175 39287
rect 16117 39247 16175 39253
rect 17405 39287 17463 39293
rect 17405 39253 17417 39287
rect 17451 39253 17463 39287
rect 17512 39284 17540 39460
rect 17586 39448 17592 39500
rect 17644 39488 17650 39500
rect 17957 39491 18015 39497
rect 17957 39488 17969 39491
rect 17644 39460 17969 39488
rect 17644 39448 17650 39460
rect 17957 39457 17969 39460
rect 18003 39457 18015 39491
rect 17957 39451 18015 39457
rect 18046 39448 18052 39500
rect 18104 39448 18110 39500
rect 20165 39491 20223 39497
rect 20165 39457 20177 39491
rect 20211 39488 20223 39491
rect 20346 39488 20352 39500
rect 20211 39460 20352 39488
rect 20211 39457 20223 39460
rect 20165 39451 20223 39457
rect 20346 39448 20352 39460
rect 20404 39448 20410 39500
rect 21082 39448 21088 39500
rect 21140 39488 21146 39500
rect 21269 39491 21327 39497
rect 21269 39488 21281 39491
rect 21140 39460 21281 39488
rect 21140 39448 21146 39460
rect 21269 39457 21281 39460
rect 21315 39457 21327 39491
rect 21269 39451 21327 39457
rect 21634 39448 21640 39500
rect 21692 39488 21698 39500
rect 22373 39491 22431 39497
rect 22373 39488 22385 39491
rect 21692 39460 22385 39488
rect 21692 39448 21698 39460
rect 22373 39457 22385 39460
rect 22419 39457 22431 39491
rect 22373 39451 22431 39457
rect 22465 39491 22523 39497
rect 22465 39457 22477 39491
rect 22511 39488 22523 39491
rect 22830 39488 22836 39500
rect 22511 39460 22836 39488
rect 22511 39457 22523 39460
rect 22465 39451 22523 39457
rect 17865 39423 17923 39429
rect 17865 39389 17877 39423
rect 17911 39420 17923 39423
rect 18064 39420 18092 39448
rect 21177 39423 21235 39429
rect 21177 39420 21189 39423
rect 17911 39392 18092 39420
rect 19306 39392 21189 39420
rect 17911 39389 17923 39392
rect 17865 39383 17923 39389
rect 17586 39312 17592 39364
rect 17644 39352 17650 39364
rect 17773 39355 17831 39361
rect 17773 39352 17785 39355
rect 17644 39324 17785 39352
rect 17644 39312 17650 39324
rect 17773 39321 17785 39324
rect 17819 39321 17831 39355
rect 17773 39315 17831 39321
rect 17954 39312 17960 39364
rect 18012 39352 18018 39364
rect 19306 39352 19334 39392
rect 21177 39389 21189 39392
rect 21223 39420 21235 39423
rect 21223 39392 22094 39420
rect 21223 39389 21235 39392
rect 21177 39383 21235 39389
rect 18012 39324 19334 39352
rect 18012 39312 18018 39324
rect 19610 39312 19616 39364
rect 19668 39352 19674 39364
rect 21085 39355 21143 39361
rect 19668 39324 20024 39352
rect 19668 39312 19674 39324
rect 18966 39284 18972 39296
rect 17512 39256 18972 39284
rect 17405 39247 17463 39253
rect 18966 39244 18972 39256
rect 19024 39244 19030 39296
rect 19886 39244 19892 39296
rect 19944 39244 19950 39296
rect 19996 39293 20024 39324
rect 21085 39321 21097 39355
rect 21131 39352 21143 39355
rect 21818 39352 21824 39364
rect 21131 39324 21824 39352
rect 21131 39321 21143 39324
rect 21085 39315 21143 39321
rect 21818 39312 21824 39324
rect 21876 39312 21882 39364
rect 22066 39352 22094 39392
rect 22186 39380 22192 39432
rect 22244 39420 22250 39432
rect 22480 39420 22508 39451
rect 22830 39448 22836 39460
rect 22888 39448 22894 39500
rect 25038 39448 25044 39500
rect 25096 39488 25102 39500
rect 25133 39491 25191 39497
rect 25133 39488 25145 39491
rect 25096 39460 25145 39488
rect 25096 39448 25102 39460
rect 25133 39457 25145 39460
rect 25179 39457 25191 39491
rect 25133 39451 25191 39457
rect 22244 39392 22508 39420
rect 22244 39380 22250 39392
rect 24026 39380 24032 39432
rect 24084 39380 24090 39432
rect 24946 39380 24952 39432
rect 25004 39380 25010 39432
rect 22462 39352 22468 39364
rect 22066 39324 22468 39352
rect 22462 39312 22468 39324
rect 22520 39352 22526 39364
rect 25406 39352 25412 39364
rect 22520 39324 25412 39352
rect 22520 39312 22526 39324
rect 25406 39312 25412 39324
rect 25464 39312 25470 39364
rect 19981 39287 20039 39293
rect 19981 39253 19993 39287
rect 20027 39284 20039 39287
rect 20622 39284 20628 39296
rect 20027 39256 20628 39284
rect 20027 39253 20039 39256
rect 19981 39247 20039 39253
rect 20622 39244 20628 39256
rect 20680 39244 20686 39296
rect 21910 39244 21916 39296
rect 21968 39244 21974 39296
rect 22278 39244 22284 39296
rect 22336 39244 22342 39296
rect 23845 39287 23903 39293
rect 23845 39253 23857 39287
rect 23891 39284 23903 39287
rect 24302 39284 24308 39296
rect 23891 39256 24308 39284
rect 23891 39253 23903 39256
rect 23845 39247 23903 39253
rect 24302 39244 24308 39256
rect 24360 39244 24366 39296
rect 25038 39244 25044 39296
rect 25096 39244 25102 39296
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 9677 39083 9735 39089
rect 9677 39049 9689 39083
rect 9723 39080 9735 39083
rect 9766 39080 9772 39092
rect 9723 39052 9772 39080
rect 9723 39049 9735 39052
rect 9677 39043 9735 39049
rect 9766 39040 9772 39052
rect 9824 39040 9830 39092
rect 11793 39083 11851 39089
rect 11793 39049 11805 39083
rect 11839 39080 11851 39083
rect 11882 39080 11888 39092
rect 11839 39052 11888 39080
rect 11839 39049 11851 39052
rect 11793 39043 11851 39049
rect 11882 39040 11888 39052
rect 11940 39040 11946 39092
rect 13998 39040 14004 39092
rect 14056 39040 14062 39092
rect 15933 39083 15991 39089
rect 15933 39049 15945 39083
rect 15979 39080 15991 39083
rect 16850 39080 16856 39092
rect 15979 39052 16856 39080
rect 15979 39049 15991 39052
rect 15933 39043 15991 39049
rect 16850 39040 16856 39052
rect 16908 39040 16914 39092
rect 18598 39080 18604 39092
rect 17972 39052 18604 39080
rect 10137 39015 10195 39021
rect 10137 38981 10149 39015
rect 10183 39012 10195 39015
rect 12710 39012 12716 39024
rect 10183 38984 12716 39012
rect 10183 38981 10195 38984
rect 10137 38975 10195 38981
rect 12710 38972 12716 38984
rect 12768 38972 12774 39024
rect 12986 38972 12992 39024
rect 13044 39012 13050 39024
rect 16574 39012 16580 39024
rect 13044 38984 16580 39012
rect 13044 38972 13050 38984
rect 16574 38972 16580 38984
rect 16632 39012 16638 39024
rect 17310 39012 17316 39024
rect 16632 38984 17316 39012
rect 16632 38972 16638 38984
rect 17310 38972 17316 38984
rect 17368 38972 17374 39024
rect 17972 39021 18000 39052
rect 18598 39040 18604 39052
rect 18656 39080 18662 39092
rect 18656 39052 19288 39080
rect 18656 39040 18662 39052
rect 17957 39015 18015 39021
rect 17957 38981 17969 39015
rect 18003 38981 18015 39015
rect 17957 38975 18015 38981
rect 18414 38972 18420 39024
rect 18472 38972 18478 39024
rect 19260 39012 19288 39052
rect 19702 39040 19708 39092
rect 19760 39080 19766 39092
rect 20349 39083 20407 39089
rect 20349 39080 20361 39083
rect 19760 39052 20361 39080
rect 19760 39040 19766 39052
rect 20349 39049 20361 39052
rect 20395 39049 20407 39083
rect 20349 39043 20407 39049
rect 22370 39040 22376 39092
rect 22428 39080 22434 39092
rect 22465 39083 22523 39089
rect 22465 39080 22477 39083
rect 22428 39052 22477 39080
rect 22428 39040 22434 39052
rect 22465 39049 22477 39052
rect 22511 39049 22523 39083
rect 25133 39083 25191 39089
rect 25133 39080 25145 39083
rect 22465 39043 22523 39049
rect 23308 39052 25145 39080
rect 19260 38984 20392 39012
rect 934 38904 940 38956
rect 992 38944 998 38956
rect 1765 38947 1823 38953
rect 1765 38944 1777 38947
rect 992 38916 1777 38944
rect 992 38904 998 38916
rect 1765 38913 1777 38916
rect 1811 38913 1823 38947
rect 1765 38907 1823 38913
rect 10042 38904 10048 38956
rect 10100 38904 10106 38956
rect 12161 38947 12219 38953
rect 12161 38913 12173 38947
rect 12207 38944 12219 38947
rect 13173 38947 13231 38953
rect 13173 38944 13185 38947
rect 12207 38916 13185 38944
rect 12207 38913 12219 38916
rect 12161 38907 12219 38913
rect 13173 38913 13185 38916
rect 13219 38913 13231 38947
rect 13173 38907 13231 38913
rect 15838 38904 15844 38956
rect 15896 38904 15902 38956
rect 20257 38947 20315 38953
rect 20257 38913 20269 38947
rect 20303 38913 20315 38947
rect 20364 38944 20392 38984
rect 21082 38972 21088 39024
rect 21140 39012 21146 39024
rect 22738 39012 22744 39024
rect 21140 38984 22744 39012
rect 21140 38972 21146 38984
rect 22738 38972 22744 38984
rect 22796 39012 22802 39024
rect 23308 39012 23336 39052
rect 25133 39049 25145 39052
rect 25179 39049 25191 39083
rect 25133 39043 25191 39049
rect 22796 38984 23336 39012
rect 22796 38972 22802 38984
rect 24394 38972 24400 39024
rect 24452 38972 24458 39024
rect 22373 38947 22431 38953
rect 20364 38916 22094 38944
rect 20257 38907 20315 38913
rect 9306 38836 9312 38888
rect 9364 38876 9370 38888
rect 10229 38879 10287 38885
rect 10229 38876 10241 38879
rect 9364 38848 10241 38876
rect 9364 38836 9370 38848
rect 10229 38845 10241 38848
rect 10275 38845 10287 38879
rect 10229 38839 10287 38845
rect 12250 38836 12256 38888
rect 12308 38836 12314 38888
rect 12345 38879 12403 38885
rect 12345 38845 12357 38879
rect 12391 38845 12403 38879
rect 12345 38839 12403 38845
rect 9490 38768 9496 38820
rect 9548 38808 9554 38820
rect 9548 38780 11284 38808
rect 9548 38768 9554 38780
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38740 1639 38743
rect 1854 38740 1860 38752
rect 1627 38712 1860 38740
rect 1627 38709 1639 38712
rect 1581 38703 1639 38709
rect 1854 38700 1860 38712
rect 1912 38700 1918 38752
rect 8662 38700 8668 38752
rect 8720 38700 8726 38752
rect 11057 38743 11115 38749
rect 11057 38709 11069 38743
rect 11103 38740 11115 38743
rect 11146 38740 11152 38752
rect 11103 38712 11152 38740
rect 11103 38709 11115 38712
rect 11057 38703 11115 38709
rect 11146 38700 11152 38712
rect 11204 38700 11210 38752
rect 11256 38740 11284 38780
rect 11606 38768 11612 38820
rect 11664 38808 11670 38820
rect 12360 38808 12388 38839
rect 13814 38836 13820 38888
rect 13872 38876 13878 38888
rect 14093 38879 14151 38885
rect 14093 38876 14105 38879
rect 13872 38848 14105 38876
rect 13872 38836 13878 38848
rect 14093 38845 14105 38848
rect 14139 38845 14151 38879
rect 14093 38839 14151 38845
rect 14277 38879 14335 38885
rect 14277 38845 14289 38879
rect 14323 38876 14335 38879
rect 14550 38876 14556 38888
rect 14323 38848 14556 38876
rect 14323 38845 14335 38848
rect 14277 38839 14335 38845
rect 14550 38836 14556 38848
rect 14608 38836 14614 38888
rect 16022 38836 16028 38888
rect 16080 38836 16086 38888
rect 17034 38836 17040 38888
rect 17092 38876 17098 38888
rect 17681 38879 17739 38885
rect 17681 38876 17693 38879
rect 17092 38848 17693 38876
rect 17092 38836 17098 38848
rect 17681 38845 17693 38848
rect 17727 38845 17739 38879
rect 20272 38876 20300 38907
rect 17681 38839 17739 38845
rect 18984 38848 20300 38876
rect 11664 38780 12388 38808
rect 13633 38811 13691 38817
rect 11664 38768 11670 38780
rect 13633 38777 13645 38811
rect 13679 38808 13691 38811
rect 16206 38808 16212 38820
rect 13679 38780 16212 38808
rect 13679 38777 13691 38780
rect 13633 38771 13691 38777
rect 16206 38768 16212 38780
rect 16264 38768 16270 38820
rect 13354 38740 13360 38752
rect 11256 38712 13360 38740
rect 13354 38700 13360 38712
rect 13412 38700 13418 38752
rect 15473 38743 15531 38749
rect 15473 38709 15485 38743
rect 15519 38740 15531 38743
rect 16482 38740 16488 38752
rect 15519 38712 16488 38740
rect 15519 38709 15531 38712
rect 15473 38703 15531 38709
rect 16482 38700 16488 38712
rect 16540 38700 16546 38752
rect 16666 38700 16672 38752
rect 16724 38740 16730 38752
rect 18984 38740 19012 38848
rect 20438 38836 20444 38888
rect 20496 38836 20502 38888
rect 19429 38811 19487 38817
rect 19429 38777 19441 38811
rect 19475 38808 19487 38811
rect 19610 38808 19616 38820
rect 19475 38780 19616 38808
rect 19475 38777 19487 38780
rect 19429 38771 19487 38777
rect 19610 38768 19616 38780
rect 19668 38768 19674 38820
rect 22066 38808 22094 38916
rect 22373 38913 22385 38947
rect 22419 38944 22431 38947
rect 22830 38944 22836 38956
rect 22419 38916 22836 38944
rect 22419 38913 22431 38916
rect 22373 38907 22431 38913
rect 22830 38904 22836 38916
rect 22888 38904 22894 38956
rect 22557 38879 22615 38885
rect 22557 38845 22569 38879
rect 22603 38845 22615 38879
rect 22557 38839 22615 38845
rect 22572 38808 22600 38839
rect 23382 38836 23388 38888
rect 23440 38836 23446 38888
rect 23661 38879 23719 38885
rect 23661 38845 23673 38879
rect 23707 38876 23719 38879
rect 24210 38876 24216 38888
rect 23707 38848 24216 38876
rect 23707 38845 23719 38848
rect 23661 38839 23719 38845
rect 24210 38836 24216 38848
rect 24268 38836 24274 38888
rect 22066 38780 22600 38808
rect 16724 38712 19012 38740
rect 16724 38700 16730 38712
rect 19518 38700 19524 38752
rect 19576 38740 19582 38752
rect 19889 38743 19947 38749
rect 19889 38740 19901 38743
rect 19576 38712 19901 38740
rect 19576 38700 19582 38712
rect 19889 38709 19901 38712
rect 19935 38709 19947 38743
rect 19889 38703 19947 38709
rect 22002 38700 22008 38752
rect 22060 38700 22066 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 6549 38539 6607 38545
rect 6549 38505 6561 38539
rect 6595 38536 6607 38539
rect 6914 38536 6920 38548
rect 6595 38508 6920 38536
rect 6595 38505 6607 38508
rect 6549 38499 6607 38505
rect 6914 38496 6920 38508
rect 6972 38496 6978 38548
rect 7558 38496 7564 38548
rect 7616 38496 7622 38548
rect 7834 38496 7840 38548
rect 7892 38496 7898 38548
rect 9398 38496 9404 38548
rect 9456 38536 9462 38548
rect 9493 38539 9551 38545
rect 9493 38536 9505 38539
rect 9456 38508 9505 38536
rect 9456 38496 9462 38508
rect 9493 38505 9505 38508
rect 9539 38505 9551 38539
rect 10689 38539 10747 38545
rect 9493 38499 9551 38505
rect 9600 38508 10088 38536
rect 7576 38468 7604 38496
rect 9600 38468 9628 38508
rect 7576 38440 9628 38468
rect 10060 38468 10088 38508
rect 10689 38505 10701 38539
rect 10735 38536 10747 38539
rect 11514 38536 11520 38548
rect 10735 38508 11520 38536
rect 10735 38505 10747 38508
rect 10689 38499 10747 38505
rect 11514 38496 11520 38508
rect 11572 38496 11578 38548
rect 11716 38508 14872 38536
rect 11238 38468 11244 38480
rect 10060 38440 11244 38468
rect 4801 38403 4859 38409
rect 4801 38369 4813 38403
rect 4847 38400 4859 38403
rect 6270 38400 6276 38412
rect 4847 38372 6276 38400
rect 4847 38369 4859 38372
rect 4801 38363 4859 38369
rect 6270 38360 6276 38372
rect 6328 38400 6334 38412
rect 7558 38400 7564 38412
rect 6328 38372 7564 38400
rect 6328 38360 6334 38372
rect 7558 38360 7564 38372
rect 7616 38360 7622 38412
rect 8496 38409 8524 38440
rect 11238 38428 11244 38440
rect 11296 38428 11302 38480
rect 11716 38468 11744 38508
rect 11348 38440 11744 38468
rect 11977 38471 12035 38477
rect 11348 38412 11376 38440
rect 11977 38437 11989 38471
rect 12023 38437 12035 38471
rect 11977 38431 12035 38437
rect 8481 38403 8539 38409
rect 8481 38369 8493 38403
rect 8527 38369 8539 38403
rect 10045 38403 10103 38409
rect 10045 38400 10057 38403
rect 8481 38363 8539 38369
rect 8772 38372 10057 38400
rect 7374 38292 7380 38344
rect 7432 38332 7438 38344
rect 8018 38332 8024 38344
rect 7432 38304 8024 38332
rect 7432 38292 7438 38304
rect 8018 38292 8024 38304
rect 8076 38292 8082 38344
rect 8205 38335 8263 38341
rect 8205 38301 8217 38335
rect 8251 38332 8263 38335
rect 8662 38332 8668 38344
rect 8251 38304 8668 38332
rect 8251 38301 8263 38304
rect 8205 38295 8263 38301
rect 8662 38292 8668 38304
rect 8720 38292 8726 38344
rect 5077 38267 5135 38273
rect 5077 38233 5089 38267
rect 5123 38233 5135 38267
rect 5077 38227 5135 38233
rect 5092 38196 5120 38227
rect 5534 38224 5540 38276
rect 5592 38224 5598 38276
rect 8772 38264 8800 38372
rect 10045 38369 10057 38372
rect 10091 38369 10103 38403
rect 10045 38363 10103 38369
rect 10318 38360 10324 38412
rect 10376 38400 10382 38412
rect 11149 38403 11207 38409
rect 11149 38400 11161 38403
rect 10376 38372 11161 38400
rect 10376 38360 10382 38372
rect 11149 38369 11161 38372
rect 11195 38369 11207 38403
rect 11149 38363 11207 38369
rect 11330 38360 11336 38412
rect 11388 38360 11394 38412
rect 9582 38292 9588 38344
rect 9640 38332 9646 38344
rect 11992 38332 12020 38431
rect 12158 38428 12164 38480
rect 12216 38468 12222 38480
rect 14844 38468 14872 38508
rect 16758 38496 16764 38548
rect 16816 38496 16822 38548
rect 20625 38539 20683 38545
rect 20625 38505 20637 38539
rect 20671 38536 20683 38539
rect 22278 38536 22284 38548
rect 20671 38508 22284 38536
rect 20671 38505 20683 38508
rect 20625 38499 20683 38505
rect 22278 38496 22284 38508
rect 22336 38496 22342 38548
rect 22554 38496 22560 38548
rect 22612 38536 22618 38548
rect 23474 38536 23480 38548
rect 22612 38508 23480 38536
rect 22612 38496 22618 38508
rect 23474 38496 23480 38508
rect 23532 38496 23538 38548
rect 21821 38471 21879 38477
rect 12216 38440 13308 38468
rect 14844 38440 17356 38468
rect 12216 38428 12222 38440
rect 12342 38360 12348 38412
rect 12400 38400 12406 38412
rect 12437 38403 12495 38409
rect 12437 38400 12449 38403
rect 12400 38372 12449 38400
rect 12400 38360 12406 38372
rect 12437 38369 12449 38372
rect 12483 38369 12495 38403
rect 12437 38363 12495 38369
rect 12529 38403 12587 38409
rect 12529 38369 12541 38403
rect 12575 38369 12587 38403
rect 12529 38363 12587 38369
rect 12544 38332 12572 38363
rect 9640 38304 12020 38332
rect 12406 38304 12572 38332
rect 13280 38332 13308 38440
rect 13354 38360 13360 38412
rect 13412 38400 13418 38412
rect 14829 38403 14887 38409
rect 14829 38400 14841 38403
rect 13412 38372 14841 38400
rect 13412 38360 13418 38372
rect 14829 38369 14841 38372
rect 14875 38369 14887 38403
rect 14829 38363 14887 38369
rect 14921 38403 14979 38409
rect 14921 38369 14933 38403
rect 14967 38369 14979 38403
rect 14921 38363 14979 38369
rect 14550 38332 14556 38344
rect 13280 38304 14556 38332
rect 9640 38292 9646 38304
rect 7852 38236 8800 38264
rect 7852 38208 7880 38236
rect 9766 38224 9772 38276
rect 9824 38264 9830 38276
rect 9953 38267 10011 38273
rect 9953 38264 9965 38267
rect 9824 38236 9965 38264
rect 9824 38224 9830 38236
rect 9953 38233 9965 38236
rect 9999 38233 10011 38267
rect 11330 38264 11336 38276
rect 9953 38227 10011 38233
rect 10060 38236 11336 38264
rect 7834 38196 7840 38208
rect 5092 38168 7840 38196
rect 7834 38156 7840 38168
rect 7892 38156 7898 38208
rect 8018 38156 8024 38208
rect 8076 38196 8082 38208
rect 8297 38199 8355 38205
rect 8297 38196 8309 38199
rect 8076 38168 8309 38196
rect 8076 38156 8082 38168
rect 8297 38165 8309 38168
rect 8343 38196 8355 38199
rect 8386 38196 8392 38208
rect 8343 38168 8392 38196
rect 8343 38165 8355 38168
rect 8297 38159 8355 38165
rect 8386 38156 8392 38168
rect 8444 38156 8450 38208
rect 9861 38199 9919 38205
rect 9861 38165 9873 38199
rect 9907 38196 9919 38199
rect 10060 38196 10088 38236
rect 11330 38224 11336 38236
rect 11388 38224 11394 38276
rect 12406 38264 12434 38304
rect 14550 38292 14556 38304
rect 14608 38332 14614 38344
rect 14936 38332 14964 38363
rect 16298 38360 16304 38412
rect 16356 38360 16362 38412
rect 17218 38360 17224 38412
rect 17276 38360 17282 38412
rect 17328 38409 17356 38440
rect 21821 38437 21833 38471
rect 21867 38468 21879 38471
rect 22094 38468 22100 38480
rect 21867 38440 22100 38468
rect 21867 38437 21879 38440
rect 21821 38431 21879 38437
rect 22094 38428 22100 38440
rect 22152 38428 22158 38480
rect 25682 38468 25688 38480
rect 22296 38440 25688 38468
rect 17313 38403 17371 38409
rect 17313 38369 17325 38403
rect 17359 38369 17371 38403
rect 17313 38363 17371 38369
rect 19334 38360 19340 38412
rect 19392 38400 19398 38412
rect 19889 38403 19947 38409
rect 19889 38400 19901 38403
rect 19392 38372 19901 38400
rect 19392 38360 19398 38372
rect 19889 38369 19901 38372
rect 19935 38369 19947 38403
rect 19889 38363 19947 38369
rect 20070 38360 20076 38412
rect 20128 38360 20134 38412
rect 21266 38360 21272 38412
rect 21324 38360 21330 38412
rect 22296 38400 22324 38440
rect 25682 38428 25688 38440
rect 25740 38428 25746 38480
rect 21376 38372 22324 38400
rect 22465 38403 22523 38409
rect 21376 38332 21404 38372
rect 22465 38369 22477 38403
rect 22511 38400 22523 38403
rect 22554 38400 22560 38412
rect 22511 38372 22560 38400
rect 22511 38369 22523 38372
rect 22465 38363 22523 38369
rect 22554 38360 22560 38372
rect 22612 38360 22618 38412
rect 23290 38360 23296 38412
rect 23348 38400 23354 38412
rect 23569 38403 23627 38409
rect 23569 38400 23581 38403
rect 23348 38372 23581 38400
rect 23348 38360 23354 38372
rect 23569 38369 23581 38372
rect 23615 38369 23627 38403
rect 23569 38363 23627 38369
rect 14608 38304 14964 38332
rect 21008 38304 21404 38332
rect 14608 38292 14614 38304
rect 11992 38236 12434 38264
rect 14737 38267 14795 38273
rect 9907 38168 10088 38196
rect 9907 38165 9919 38168
rect 9861 38159 9919 38165
rect 11054 38156 11060 38208
rect 11112 38156 11118 38208
rect 11238 38156 11244 38208
rect 11296 38196 11302 38208
rect 11992 38196 12020 38236
rect 14737 38233 14749 38267
rect 14783 38264 14795 38267
rect 17586 38264 17592 38276
rect 14783 38236 15700 38264
rect 14783 38233 14795 38236
rect 14737 38227 14795 38233
rect 15672 38208 15700 38236
rect 15764 38236 17592 38264
rect 11296 38168 12020 38196
rect 11296 38156 11302 38168
rect 12342 38156 12348 38208
rect 12400 38156 12406 38208
rect 14366 38156 14372 38208
rect 14424 38156 14430 38208
rect 15654 38156 15660 38208
rect 15712 38156 15718 38208
rect 15764 38205 15792 38236
rect 17586 38224 17592 38236
rect 17644 38224 17650 38276
rect 18598 38224 18604 38276
rect 18656 38264 18662 38276
rect 19797 38267 19855 38273
rect 19797 38264 19809 38267
rect 18656 38236 19809 38264
rect 18656 38224 18662 38236
rect 19797 38233 19809 38236
rect 19843 38233 19855 38267
rect 19797 38227 19855 38233
rect 19978 38224 19984 38276
rect 20036 38264 20042 38276
rect 21008 38273 21036 38304
rect 21542 38292 21548 38344
rect 21600 38332 21606 38344
rect 23477 38335 23535 38341
rect 23477 38332 23489 38335
rect 21600 38304 23489 38332
rect 21600 38292 21606 38304
rect 23477 38301 23489 38304
rect 23523 38301 23535 38335
rect 23477 38295 23535 38301
rect 25317 38335 25375 38341
rect 25317 38301 25329 38335
rect 25363 38332 25375 38335
rect 25406 38332 25412 38344
rect 25363 38304 25412 38332
rect 25363 38301 25375 38304
rect 25317 38295 25375 38301
rect 25406 38292 25412 38304
rect 25464 38292 25470 38344
rect 20993 38267 21051 38273
rect 20993 38264 21005 38267
rect 20036 38236 21005 38264
rect 20036 38224 20042 38236
rect 20993 38233 21005 38236
rect 21039 38233 21051 38267
rect 20993 38227 21051 38233
rect 21450 38224 21456 38276
rect 21508 38264 21514 38276
rect 23385 38267 23443 38273
rect 23385 38264 23397 38267
rect 21508 38236 23397 38264
rect 21508 38224 21514 38236
rect 23385 38233 23397 38236
rect 23431 38233 23443 38267
rect 23385 38227 23443 38233
rect 15749 38199 15807 38205
rect 15749 38165 15761 38199
rect 15795 38165 15807 38199
rect 15749 38159 15807 38165
rect 16114 38156 16120 38208
rect 16172 38156 16178 38208
rect 16206 38156 16212 38208
rect 16264 38156 16270 38208
rect 17126 38156 17132 38208
rect 17184 38156 17190 38208
rect 19429 38199 19487 38205
rect 19429 38165 19441 38199
rect 19475 38196 19487 38199
rect 20254 38196 20260 38208
rect 19475 38168 20260 38196
rect 19475 38165 19487 38168
rect 19429 38159 19487 38165
rect 20254 38156 20260 38168
rect 20312 38156 20318 38208
rect 20714 38156 20720 38208
rect 20772 38196 20778 38208
rect 21085 38199 21143 38205
rect 21085 38196 21097 38199
rect 20772 38168 21097 38196
rect 20772 38156 20778 38168
rect 21085 38165 21097 38168
rect 21131 38165 21143 38199
rect 21085 38159 21143 38165
rect 21818 38156 21824 38208
rect 21876 38196 21882 38208
rect 22189 38199 22247 38205
rect 22189 38196 22201 38199
rect 21876 38168 22201 38196
rect 21876 38156 21882 38168
rect 22189 38165 22201 38168
rect 22235 38165 22247 38199
rect 22189 38159 22247 38165
rect 22281 38199 22339 38205
rect 22281 38165 22293 38199
rect 22327 38196 22339 38199
rect 22462 38196 22468 38208
rect 22327 38168 22468 38196
rect 22327 38165 22339 38168
rect 22281 38159 22339 38165
rect 22462 38156 22468 38168
rect 22520 38156 22526 38208
rect 23017 38199 23075 38205
rect 23017 38165 23029 38199
rect 23063 38196 23075 38199
rect 23658 38196 23664 38208
rect 23063 38168 23664 38196
rect 23063 38165 23075 38168
rect 23017 38159 23075 38165
rect 23658 38156 23664 38168
rect 23716 38156 23722 38208
rect 25130 38156 25136 38208
rect 25188 38156 25194 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5997 37995 6055 38001
rect 5997 37961 6009 37995
rect 6043 37992 6055 37995
rect 6546 37992 6552 38004
rect 6043 37964 6552 37992
rect 6043 37961 6055 37964
rect 5997 37955 6055 37961
rect 6546 37952 6552 37964
rect 6604 37952 6610 38004
rect 7006 37952 7012 38004
rect 7064 37992 7070 38004
rect 10318 37992 10324 38004
rect 7064 37964 10324 37992
rect 7064 37952 7070 37964
rect 10318 37952 10324 37964
rect 10376 37952 10382 38004
rect 10505 37995 10563 38001
rect 10505 37961 10517 37995
rect 10551 37992 10563 37995
rect 11146 37992 11152 38004
rect 10551 37964 11152 37992
rect 10551 37961 10563 37964
rect 10505 37955 10563 37961
rect 11146 37952 11152 37964
rect 11204 37952 11210 38004
rect 11330 37952 11336 38004
rect 11388 37992 11394 38004
rect 12802 37992 12808 38004
rect 11388 37964 12808 37992
rect 11388 37952 11394 37964
rect 12802 37952 12808 37964
rect 12860 37952 12866 38004
rect 12897 37995 12955 38001
rect 12897 37961 12909 37995
rect 12943 37992 12955 37995
rect 15838 37992 15844 38004
rect 12943 37964 15844 37992
rect 12943 37961 12955 37964
rect 12897 37955 12955 37961
rect 15838 37952 15844 37964
rect 15896 37952 15902 38004
rect 17328 37964 18736 37992
rect 5534 37884 5540 37936
rect 5592 37884 5598 37936
rect 8294 37884 8300 37936
rect 8352 37884 8358 37936
rect 10336 37924 10364 37952
rect 13357 37927 13415 37933
rect 13357 37924 13369 37927
rect 10336 37896 13369 37924
rect 13357 37893 13369 37896
rect 13403 37893 13415 37927
rect 13357 37887 13415 37893
rect 14182 37884 14188 37936
rect 14240 37924 14246 37936
rect 15381 37927 15439 37933
rect 15381 37924 15393 37927
rect 14240 37896 15393 37924
rect 14240 37884 14246 37896
rect 15381 37893 15393 37896
rect 15427 37893 15439 37927
rect 15381 37887 15439 37893
rect 16574 37884 16580 37936
rect 16632 37924 16638 37936
rect 17328 37933 17356 37964
rect 17313 37927 17371 37933
rect 17313 37924 17325 37927
rect 16632 37896 17325 37924
rect 16632 37884 16638 37896
rect 17313 37893 17325 37896
rect 17359 37893 17371 37927
rect 18708 37924 18736 37964
rect 18782 37952 18788 38004
rect 18840 37952 18846 38004
rect 19610 37992 19616 38004
rect 19352 37964 19616 37992
rect 19352 37924 19380 37964
rect 19610 37952 19616 37964
rect 19668 37952 19674 38004
rect 20533 37995 20591 38001
rect 20533 37961 20545 37995
rect 20579 37992 20591 37995
rect 22370 37992 22376 38004
rect 20579 37964 22376 37992
rect 20579 37961 20591 37964
rect 20533 37955 20591 37961
rect 22370 37952 22376 37964
rect 22428 37952 22434 38004
rect 22738 37952 22744 38004
rect 22796 37992 22802 38004
rect 23750 37992 23756 38004
rect 22796 37964 23756 37992
rect 22796 37952 22802 37964
rect 23750 37952 23756 37964
rect 23808 37952 23814 38004
rect 24210 37952 24216 38004
rect 24268 37992 24274 38004
rect 25317 37995 25375 38001
rect 25317 37992 25329 37995
rect 24268 37964 25329 37992
rect 24268 37952 24274 37964
rect 25317 37961 25329 37964
rect 25363 37961 25375 37995
rect 25317 37955 25375 37961
rect 18708 37896 19380 37924
rect 17313 37887 17371 37893
rect 19426 37884 19432 37936
rect 19484 37924 19490 37936
rect 22005 37927 22063 37933
rect 22005 37924 22017 37927
rect 19484 37896 22017 37924
rect 19484 37884 19490 37896
rect 22005 37893 22017 37896
rect 22051 37893 22063 37927
rect 22005 37887 22063 37893
rect 23290 37884 23296 37936
rect 23348 37924 23354 37936
rect 23845 37927 23903 37933
rect 23845 37924 23857 37927
rect 23348 37896 23857 37924
rect 23348 37884 23354 37896
rect 23845 37893 23857 37896
rect 23891 37893 23903 37927
rect 23845 37887 23903 37893
rect 24486 37884 24492 37936
rect 24544 37884 24550 37936
rect 7558 37816 7564 37868
rect 7616 37816 7622 37868
rect 10226 37816 10232 37868
rect 10284 37856 10290 37868
rect 10284 37828 10732 37856
rect 10284 37816 10290 37828
rect 10704 37800 10732 37828
rect 11054 37816 11060 37868
rect 11112 37856 11118 37868
rect 11885 37859 11943 37865
rect 11885 37856 11897 37859
rect 11112 37828 11897 37856
rect 11112 37816 11118 37828
rect 11885 37825 11897 37828
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 13265 37859 13323 37865
rect 13265 37825 13277 37859
rect 13311 37856 13323 37859
rect 14277 37859 14335 37865
rect 14277 37856 14289 37859
rect 13311 37828 14289 37856
rect 13311 37825 13323 37828
rect 13265 37819 13323 37825
rect 14277 37825 14289 37828
rect 14323 37825 14335 37859
rect 14277 37819 14335 37825
rect 15286 37816 15292 37868
rect 15344 37816 15350 37868
rect 16114 37816 16120 37868
rect 16172 37856 16178 37868
rect 16301 37859 16359 37865
rect 16301 37856 16313 37859
rect 16172 37828 16313 37856
rect 16172 37816 16178 37828
rect 16301 37825 16313 37828
rect 16347 37825 16359 37859
rect 16301 37819 16359 37825
rect 18414 37816 18420 37868
rect 18472 37856 18478 37868
rect 19058 37856 19064 37868
rect 18472 37828 19064 37856
rect 18472 37816 18478 37828
rect 19058 37816 19064 37828
rect 19116 37816 19122 37868
rect 4249 37791 4307 37797
rect 4249 37757 4261 37791
rect 4295 37757 4307 37791
rect 4249 37751 4307 37757
rect 4264 37652 4292 37751
rect 4522 37748 4528 37800
rect 4580 37748 4586 37800
rect 7837 37791 7895 37797
rect 7837 37757 7849 37791
rect 7883 37788 7895 37791
rect 9306 37788 9312 37800
rect 7883 37760 9312 37788
rect 7883 37757 7895 37760
rect 7837 37751 7895 37757
rect 9306 37748 9312 37760
rect 9364 37748 9370 37800
rect 9585 37791 9643 37797
rect 9585 37757 9597 37791
rect 9631 37757 9643 37791
rect 9585 37751 9643 37757
rect 9030 37680 9036 37732
rect 9088 37720 9094 37732
rect 9600 37720 9628 37751
rect 10594 37748 10600 37800
rect 10652 37748 10658 37800
rect 10686 37748 10692 37800
rect 10744 37748 10750 37800
rect 11514 37748 11520 37800
rect 11572 37788 11578 37800
rect 13541 37791 13599 37797
rect 11572 37760 12434 37788
rect 11572 37748 11578 37760
rect 9088 37692 9628 37720
rect 10137 37723 10195 37729
rect 9088 37680 9094 37692
rect 10137 37689 10149 37723
rect 10183 37720 10195 37723
rect 12066 37720 12072 37732
rect 10183 37692 12072 37720
rect 10183 37689 10195 37692
rect 10137 37683 10195 37689
rect 12066 37680 12072 37692
rect 12124 37680 12130 37732
rect 12406 37720 12434 37760
rect 13541 37757 13553 37791
rect 13587 37788 13599 37791
rect 14182 37788 14188 37800
rect 13587 37760 14188 37788
rect 13587 37757 13599 37760
rect 13541 37751 13599 37757
rect 14182 37748 14188 37760
rect 14240 37748 14246 37800
rect 14918 37748 14924 37800
rect 14976 37788 14982 37800
rect 15473 37791 15531 37797
rect 15473 37788 15485 37791
rect 14976 37760 15485 37788
rect 14976 37748 14982 37760
rect 15473 37757 15485 37760
rect 15519 37757 15531 37791
rect 15473 37751 15531 37757
rect 17034 37748 17040 37800
rect 17092 37748 17098 37800
rect 17862 37748 17868 37800
rect 17920 37788 17926 37800
rect 20625 37791 20683 37797
rect 20625 37788 20637 37791
rect 17920 37760 20637 37788
rect 17920 37748 17926 37760
rect 20625 37757 20637 37760
rect 20671 37757 20683 37791
rect 20625 37751 20683 37757
rect 20717 37791 20775 37797
rect 20717 37757 20729 37791
rect 20763 37757 20775 37791
rect 20717 37751 20775 37757
rect 13814 37720 13820 37732
rect 12406 37692 13820 37720
rect 13814 37680 13820 37692
rect 13872 37680 13878 37732
rect 16758 37720 16764 37732
rect 14844 37692 16764 37720
rect 4982 37652 4988 37664
rect 4264 37624 4988 37652
rect 4982 37612 4988 37624
rect 5040 37612 5046 37664
rect 11054 37612 11060 37664
rect 11112 37652 11118 37664
rect 12158 37652 12164 37664
rect 11112 37624 12164 37652
rect 11112 37612 11118 37624
rect 12158 37612 12164 37624
rect 12216 37612 12222 37664
rect 12802 37612 12808 37664
rect 12860 37652 12866 37664
rect 14844 37652 14872 37692
rect 16758 37680 16764 37692
rect 16816 37680 16822 37732
rect 20530 37680 20536 37732
rect 20588 37720 20594 37732
rect 20732 37720 20760 37751
rect 22646 37748 22652 37800
rect 22704 37788 22710 37800
rect 22741 37791 22799 37797
rect 22741 37788 22753 37791
rect 22704 37760 22753 37788
rect 22704 37748 22710 37760
rect 22741 37757 22753 37760
rect 22787 37788 22799 37791
rect 23382 37788 23388 37800
rect 22787 37760 23388 37788
rect 22787 37757 22799 37760
rect 22741 37751 22799 37757
rect 23382 37748 23388 37760
rect 23440 37788 23446 37800
rect 23569 37791 23627 37797
rect 23569 37788 23581 37791
rect 23440 37760 23581 37788
rect 23440 37748 23446 37760
rect 23569 37757 23581 37760
rect 23615 37757 23627 37791
rect 23569 37751 23627 37757
rect 20588 37692 20760 37720
rect 20588 37680 20594 37692
rect 12860 37624 14872 37652
rect 12860 37612 12866 37624
rect 14918 37612 14924 37664
rect 14976 37612 14982 37664
rect 18046 37612 18052 37664
rect 18104 37652 18110 37664
rect 18506 37652 18512 37664
rect 18104 37624 18512 37652
rect 18104 37612 18110 37624
rect 18506 37612 18512 37624
rect 18564 37612 18570 37664
rect 19610 37612 19616 37664
rect 19668 37612 19674 37664
rect 20165 37655 20223 37661
rect 20165 37621 20177 37655
rect 20211 37652 20223 37655
rect 20990 37652 20996 37664
rect 20211 37624 20996 37652
rect 20211 37621 20223 37624
rect 20165 37615 20223 37621
rect 20990 37612 20996 37624
rect 21048 37612 21054 37664
rect 21542 37612 21548 37664
rect 21600 37652 21606 37664
rect 25222 37652 25228 37664
rect 21600 37624 25228 37652
rect 21600 37612 21606 37624
rect 25222 37612 25228 37624
rect 25280 37612 25286 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 6178 37408 6184 37460
rect 6236 37448 6242 37460
rect 7006 37448 7012 37460
rect 6236 37420 7012 37448
rect 6236 37408 6242 37420
rect 7006 37408 7012 37420
rect 7064 37408 7070 37460
rect 10686 37408 10692 37460
rect 10744 37448 10750 37460
rect 10744 37420 15516 37448
rect 10744 37408 10750 37420
rect 8386 37340 8392 37392
rect 8444 37380 8450 37392
rect 11514 37380 11520 37392
rect 8444 37352 11520 37380
rect 8444 37340 8450 37352
rect 11514 37340 11520 37352
rect 11572 37340 11578 37392
rect 15378 37340 15384 37392
rect 15436 37340 15442 37392
rect 15488 37380 15516 37420
rect 15654 37408 15660 37460
rect 15712 37448 15718 37460
rect 22370 37448 22376 37460
rect 15712 37420 22376 37448
rect 15712 37408 15718 37420
rect 22370 37408 22376 37420
rect 22428 37448 22434 37460
rect 22738 37448 22744 37460
rect 22428 37420 22744 37448
rect 22428 37408 22434 37420
rect 22738 37408 22744 37420
rect 22796 37408 22802 37460
rect 16390 37380 16396 37392
rect 15488 37352 16396 37380
rect 16390 37340 16396 37352
rect 16448 37340 16454 37392
rect 17218 37380 17224 37392
rect 16592 37352 17224 37380
rect 5537 37315 5595 37321
rect 5537 37281 5549 37315
rect 5583 37312 5595 37315
rect 6914 37312 6920 37324
rect 5583 37284 6920 37312
rect 5583 37281 5595 37284
rect 5537 37275 5595 37281
rect 6914 37272 6920 37284
rect 6972 37272 6978 37324
rect 7006 37272 7012 37324
rect 7064 37312 7070 37324
rect 8297 37315 8355 37321
rect 8297 37312 8309 37315
rect 7064 37284 8309 37312
rect 7064 37272 7070 37284
rect 8297 37281 8309 37284
rect 8343 37281 8355 37315
rect 8297 37275 8355 37281
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 10410 37272 10416 37324
rect 10468 37312 10474 37324
rect 11885 37315 11943 37321
rect 11885 37312 11897 37315
rect 10468 37284 11897 37312
rect 10468 37272 10474 37284
rect 11885 37281 11897 37284
rect 11931 37281 11943 37315
rect 15396 37312 15424 37340
rect 15657 37315 15715 37321
rect 15657 37312 15669 37315
rect 15396 37284 15669 37312
rect 11885 37275 11943 37281
rect 15657 37281 15669 37284
rect 15703 37312 15715 37315
rect 16206 37312 16212 37324
rect 15703 37284 16212 37312
rect 15703 37281 15715 37284
rect 15657 37275 15715 37281
rect 16206 37272 16212 37284
rect 16264 37272 16270 37324
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5040 37216 5273 37244
rect 5040 37204 5046 37216
rect 5261 37213 5273 37216
rect 5307 37213 5319 37247
rect 5261 37207 5319 37213
rect 7282 37204 7288 37256
rect 7340 37204 7346 37256
rect 8754 37204 8760 37256
rect 8812 37244 8818 37256
rect 10229 37247 10287 37253
rect 10229 37244 10241 37247
rect 8812 37216 10241 37244
rect 8812 37204 8818 37216
rect 10229 37213 10241 37216
rect 10275 37213 10287 37247
rect 13630 37244 13636 37256
rect 10229 37207 10287 37213
rect 10336 37216 13636 37244
rect 5534 37136 5540 37188
rect 5592 37176 5598 37188
rect 8113 37179 8171 37185
rect 5592 37148 6026 37176
rect 5592 37136 5598 37148
rect 8113 37145 8125 37179
rect 8159 37176 8171 37179
rect 9858 37176 9864 37188
rect 8159 37148 9864 37176
rect 8159 37145 8171 37148
rect 8113 37139 8171 37145
rect 9858 37136 9864 37148
rect 9916 37136 9922 37188
rect 7742 37068 7748 37120
rect 7800 37068 7806 37120
rect 8205 37111 8263 37117
rect 8205 37077 8217 37111
rect 8251 37108 8263 37111
rect 9769 37111 9827 37117
rect 9769 37108 9781 37111
rect 8251 37080 9781 37108
rect 8251 37077 8263 37080
rect 8205 37071 8263 37077
rect 9769 37077 9781 37080
rect 9815 37077 9827 37111
rect 9769 37071 9827 37077
rect 10134 37068 10140 37120
rect 10192 37068 10198 37120
rect 10226 37068 10232 37120
rect 10284 37108 10290 37120
rect 10336 37108 10364 37216
rect 13630 37204 13636 37216
rect 13688 37204 13694 37256
rect 15381 37247 15439 37253
rect 15381 37213 15393 37247
rect 15427 37244 15439 37247
rect 16592 37244 16620 37352
rect 17218 37340 17224 37352
rect 17276 37340 17282 37392
rect 19334 37380 19340 37392
rect 18616 37352 19340 37380
rect 17037 37315 17095 37321
rect 17037 37281 17049 37315
rect 17083 37312 17095 37315
rect 18046 37312 18052 37324
rect 17083 37284 18052 37312
rect 17083 37281 17095 37284
rect 17037 37275 17095 37281
rect 18046 37272 18052 37284
rect 18104 37272 18110 37324
rect 18616 37321 18644 37352
rect 19334 37340 19340 37352
rect 19392 37340 19398 37392
rect 18601 37315 18659 37321
rect 18156 37284 18552 37312
rect 15427 37216 16620 37244
rect 16761 37247 16819 37253
rect 15427 37213 15439 37216
rect 15381 37207 15439 37213
rect 16761 37213 16773 37247
rect 16807 37244 16819 37247
rect 18156 37244 18184 37284
rect 16807 37216 18184 37244
rect 18524 37244 18552 37284
rect 18601 37281 18613 37315
rect 18647 37281 18659 37315
rect 18601 37275 18659 37281
rect 18785 37315 18843 37321
rect 18785 37281 18797 37315
rect 18831 37312 18843 37315
rect 21082 37312 21088 37324
rect 18831 37284 21088 37312
rect 18831 37281 18843 37284
rect 18785 37275 18843 37281
rect 21082 37272 21088 37284
rect 21140 37272 21146 37324
rect 21634 37272 21640 37324
rect 21692 37312 21698 37324
rect 22186 37312 22192 37324
rect 21692 37284 22192 37312
rect 21692 37272 21698 37284
rect 22186 37272 22192 37284
rect 22244 37272 22250 37324
rect 19610 37244 19616 37256
rect 18524 37216 19616 37244
rect 16807 37213 16819 37216
rect 16761 37207 16819 37213
rect 19610 37204 19616 37216
rect 19668 37204 19674 37256
rect 21361 37247 21419 37253
rect 21361 37213 21373 37247
rect 21407 37213 21419 37247
rect 22770 37216 23704 37244
rect 21361 37207 21419 37213
rect 11701 37179 11759 37185
rect 11701 37145 11713 37179
rect 11747 37176 11759 37179
rect 15286 37176 15292 37188
rect 11747 37148 15292 37176
rect 11747 37145 11759 37148
rect 11701 37139 11759 37145
rect 15286 37136 15292 37148
rect 15344 37136 15350 37188
rect 18509 37179 18567 37185
rect 18509 37176 18521 37179
rect 17604 37148 18521 37176
rect 17604 37120 17632 37148
rect 18509 37145 18521 37148
rect 18555 37145 18567 37179
rect 18509 37139 18567 37145
rect 19426 37136 19432 37188
rect 19484 37136 19490 37188
rect 20162 37136 20168 37188
rect 20220 37136 20226 37188
rect 10284 37080 10364 37108
rect 10284 37068 10290 37080
rect 11330 37068 11336 37120
rect 11388 37068 11394 37120
rect 11793 37111 11851 37117
rect 11793 37077 11805 37111
rect 11839 37108 11851 37111
rect 15013 37111 15071 37117
rect 15013 37108 15025 37111
rect 11839 37080 15025 37108
rect 11839 37077 11851 37080
rect 11793 37071 11851 37077
rect 15013 37077 15025 37080
rect 15059 37077 15071 37111
rect 15013 37071 15071 37077
rect 15470 37068 15476 37120
rect 15528 37068 15534 37120
rect 16393 37111 16451 37117
rect 16393 37077 16405 37111
rect 16439 37108 16451 37111
rect 16666 37108 16672 37120
rect 16439 37080 16672 37108
rect 16439 37077 16451 37080
rect 16393 37071 16451 37077
rect 16666 37068 16672 37080
rect 16724 37068 16730 37120
rect 16853 37111 16911 37117
rect 16853 37077 16865 37111
rect 16899 37108 16911 37111
rect 16942 37108 16948 37120
rect 16899 37080 16948 37108
rect 16899 37077 16911 37080
rect 16853 37071 16911 37077
rect 16942 37068 16948 37080
rect 17000 37068 17006 37120
rect 17586 37068 17592 37120
rect 17644 37068 17650 37120
rect 18141 37111 18199 37117
rect 18141 37077 18153 37111
rect 18187 37108 18199 37111
rect 21174 37108 21180 37120
rect 18187 37080 21180 37108
rect 18187 37077 18199 37080
rect 18141 37071 18199 37077
rect 21174 37068 21180 37080
rect 21232 37068 21238 37120
rect 21376 37108 21404 37207
rect 22922 37136 22928 37188
rect 22980 37176 22986 37188
rect 23676 37176 23704 37216
rect 23750 37204 23756 37256
rect 23808 37204 23814 37256
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37244 24823 37247
rect 24854 37244 24860 37256
rect 24811 37216 24860 37244
rect 24811 37213 24823 37216
rect 24765 37207 24823 37213
rect 24854 37204 24860 37216
rect 24912 37204 24918 37256
rect 24486 37176 24492 37188
rect 22980 37148 23428 37176
rect 23676 37148 24492 37176
rect 22980 37136 22986 37148
rect 23400 37120 23428 37148
rect 24486 37136 24492 37148
rect 24544 37136 24550 37188
rect 22646 37108 22652 37120
rect 21376 37080 22652 37108
rect 22646 37068 22652 37080
rect 22704 37068 22710 37120
rect 23106 37068 23112 37120
rect 23164 37068 23170 37120
rect 23382 37068 23388 37120
rect 23440 37108 23446 37120
rect 23569 37111 23627 37117
rect 23569 37108 23581 37111
rect 23440 37080 23581 37108
rect 23440 37068 23446 37080
rect 23569 37077 23581 37080
rect 23615 37077 23627 37111
rect 23569 37071 23627 37077
rect 24578 37068 24584 37120
rect 24636 37068 24642 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 5166 36864 5172 36916
rect 5224 36864 5230 36916
rect 5629 36907 5687 36913
rect 5629 36873 5641 36907
rect 5675 36904 5687 36907
rect 9122 36904 9128 36916
rect 5675 36876 9128 36904
rect 5675 36873 5687 36876
rect 5629 36867 5687 36873
rect 9122 36864 9128 36876
rect 9180 36864 9186 36916
rect 9306 36864 9312 36916
rect 9364 36864 9370 36916
rect 10134 36864 10140 36916
rect 10192 36904 10198 36916
rect 10192 36876 12434 36904
rect 10192 36864 10198 36876
rect 6822 36796 6828 36848
rect 6880 36836 6886 36848
rect 8294 36836 8300 36848
rect 6880 36808 8300 36836
rect 6880 36796 6886 36808
rect 8294 36796 8300 36808
rect 8352 36796 8358 36848
rect 12406 36836 12434 36876
rect 12710 36864 12716 36916
rect 12768 36904 12774 36916
rect 12897 36907 12955 36913
rect 12897 36904 12909 36907
rect 12768 36876 12909 36904
rect 12768 36864 12774 36876
rect 12897 36873 12909 36876
rect 12943 36873 12955 36907
rect 12897 36867 12955 36873
rect 13357 36907 13415 36913
rect 13357 36873 13369 36907
rect 13403 36904 13415 36907
rect 14366 36904 14372 36916
rect 13403 36876 14372 36904
rect 13403 36873 13415 36876
rect 13357 36867 13415 36873
rect 14366 36864 14372 36876
rect 14424 36864 14430 36916
rect 15286 36864 15292 36916
rect 15344 36864 15350 36916
rect 16022 36864 16028 36916
rect 16080 36904 16086 36916
rect 16080 36876 17632 36904
rect 16080 36864 16086 36876
rect 16850 36836 16856 36848
rect 12406 36808 16856 36836
rect 16850 36796 16856 36808
rect 16908 36796 16914 36848
rect 934 36728 940 36780
rect 992 36768 998 36780
rect 1765 36771 1823 36777
rect 1765 36768 1777 36771
rect 992 36740 1777 36768
rect 992 36728 998 36740
rect 1765 36737 1777 36740
rect 1811 36737 1823 36771
rect 1765 36731 1823 36737
rect 4614 36728 4620 36780
rect 4672 36768 4678 36780
rect 5537 36771 5595 36777
rect 5537 36768 5549 36771
rect 4672 36740 5549 36768
rect 4672 36728 4678 36740
rect 5537 36737 5549 36740
rect 5583 36737 5595 36771
rect 5537 36731 5595 36737
rect 9306 36728 9312 36780
rect 9364 36768 9370 36780
rect 10137 36771 10195 36777
rect 10137 36768 10149 36771
rect 9364 36740 10149 36768
rect 9364 36728 9370 36740
rect 10137 36737 10149 36740
rect 10183 36737 10195 36771
rect 10137 36731 10195 36737
rect 13265 36771 13323 36777
rect 13265 36737 13277 36771
rect 13311 36768 13323 36771
rect 13538 36768 13544 36780
rect 13311 36740 13544 36768
rect 13311 36737 13323 36740
rect 13265 36731 13323 36737
rect 13538 36728 13544 36740
rect 13596 36728 13602 36780
rect 14829 36771 14887 36777
rect 14829 36737 14841 36771
rect 14875 36768 14887 36771
rect 15657 36771 15715 36777
rect 15657 36768 15669 36771
rect 14875 36740 15669 36768
rect 14875 36737 14887 36740
rect 14829 36731 14887 36737
rect 15657 36737 15669 36740
rect 15703 36737 15715 36771
rect 15657 36731 15715 36737
rect 15749 36771 15807 36777
rect 15749 36737 15761 36771
rect 15795 36768 15807 36771
rect 17126 36768 17132 36780
rect 15795 36740 17132 36768
rect 15795 36737 15807 36740
rect 15749 36731 15807 36737
rect 17126 36728 17132 36740
rect 17184 36768 17190 36780
rect 17494 36768 17500 36780
rect 17184 36740 17500 36768
rect 17184 36728 17190 36740
rect 17494 36728 17500 36740
rect 17552 36728 17558 36780
rect 17604 36768 17632 36876
rect 18322 36864 18328 36916
rect 18380 36904 18386 36916
rect 18417 36907 18475 36913
rect 18417 36904 18429 36907
rect 18380 36876 18429 36904
rect 18380 36864 18386 36876
rect 18417 36873 18429 36876
rect 18463 36873 18475 36907
rect 18417 36867 18475 36873
rect 19242 36864 19248 36916
rect 19300 36904 19306 36916
rect 19705 36907 19763 36913
rect 19705 36904 19717 36907
rect 19300 36876 19717 36904
rect 19300 36864 19306 36876
rect 19705 36873 19717 36876
rect 19751 36873 19763 36907
rect 19705 36867 19763 36873
rect 20165 36907 20223 36913
rect 20165 36873 20177 36907
rect 20211 36904 20223 36907
rect 22002 36904 22008 36916
rect 20211 36876 22008 36904
rect 20211 36873 20223 36876
rect 20165 36867 20223 36873
rect 22002 36864 22008 36876
rect 22060 36864 22066 36916
rect 24578 36904 24584 36916
rect 22480 36876 24584 36904
rect 17678 36796 17684 36848
rect 17736 36836 17742 36848
rect 19794 36836 19800 36848
rect 17736 36808 19800 36836
rect 17736 36796 17742 36808
rect 19794 36796 19800 36808
rect 19852 36836 19858 36848
rect 22480 36836 22508 36876
rect 24578 36864 24584 36876
rect 24636 36864 24642 36916
rect 19852 36808 22508 36836
rect 19852 36796 19858 36808
rect 22554 36796 22560 36848
rect 22612 36836 22618 36848
rect 23017 36839 23075 36845
rect 23017 36836 23029 36839
rect 22612 36808 23029 36836
rect 22612 36796 22618 36808
rect 23017 36805 23029 36808
rect 23063 36836 23075 36839
rect 23106 36836 23112 36848
rect 23063 36808 23112 36836
rect 23063 36805 23075 36808
rect 23017 36799 23075 36805
rect 23106 36796 23112 36808
rect 23164 36796 23170 36848
rect 24486 36836 24492 36848
rect 24242 36808 24492 36836
rect 24486 36796 24492 36808
rect 24544 36796 24550 36848
rect 19426 36768 19432 36780
rect 17604 36740 19432 36768
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 20073 36771 20131 36777
rect 20073 36737 20085 36771
rect 20119 36768 20131 36771
rect 22278 36768 22284 36780
rect 20119 36740 22284 36768
rect 20119 36737 20131 36740
rect 20073 36731 20131 36737
rect 22278 36728 22284 36740
rect 22336 36728 22342 36780
rect 25314 36728 25320 36780
rect 25372 36728 25378 36780
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 4522 36592 4528 36644
rect 4580 36632 4586 36644
rect 5258 36632 5264 36644
rect 4580 36604 5264 36632
rect 4580 36592 4586 36604
rect 5258 36592 5264 36604
rect 5316 36632 5322 36644
rect 5736 36632 5764 36663
rect 6086 36660 6092 36712
rect 6144 36700 6150 36712
rect 7558 36700 7564 36712
rect 6144 36672 7564 36700
rect 6144 36660 6150 36672
rect 7558 36660 7564 36672
rect 7616 36660 7622 36712
rect 7837 36703 7895 36709
rect 7837 36669 7849 36703
rect 7883 36700 7895 36703
rect 9582 36700 9588 36712
rect 7883 36672 9588 36700
rect 7883 36669 7895 36672
rect 7837 36663 7895 36669
rect 9582 36660 9588 36672
rect 9640 36660 9646 36712
rect 10226 36660 10232 36712
rect 10284 36660 10290 36712
rect 10321 36703 10379 36709
rect 10321 36669 10333 36703
rect 10367 36669 10379 36703
rect 10321 36663 10379 36669
rect 5316 36604 5764 36632
rect 5316 36592 5322 36604
rect 9490 36592 9496 36644
rect 9548 36632 9554 36644
rect 10336 36632 10364 36663
rect 13446 36660 13452 36712
rect 13504 36660 13510 36712
rect 15933 36703 15991 36709
rect 15933 36669 15945 36703
rect 15979 36700 15991 36703
rect 16206 36700 16212 36712
rect 15979 36672 16212 36700
rect 15979 36669 15991 36672
rect 15933 36663 15991 36669
rect 16206 36660 16212 36672
rect 16264 36660 16270 36712
rect 18506 36660 18512 36712
rect 18564 36660 18570 36712
rect 18601 36703 18659 36709
rect 18601 36669 18613 36703
rect 18647 36669 18659 36703
rect 18601 36663 18659 36669
rect 9548 36604 10364 36632
rect 9548 36592 9554 36604
rect 16114 36592 16120 36644
rect 16172 36632 16178 36644
rect 18049 36635 18107 36641
rect 18049 36632 18061 36635
rect 16172 36604 18061 36632
rect 16172 36592 16178 36604
rect 18049 36601 18061 36604
rect 18095 36601 18107 36635
rect 18049 36595 18107 36601
rect 18414 36592 18420 36644
rect 18472 36632 18478 36644
rect 18616 36632 18644 36663
rect 19702 36660 19708 36712
rect 19760 36700 19766 36712
rect 20257 36703 20315 36709
rect 20257 36700 20269 36703
rect 19760 36672 20269 36700
rect 19760 36660 19766 36672
rect 20257 36669 20269 36672
rect 20303 36669 20315 36703
rect 20257 36663 20315 36669
rect 22646 36660 22652 36712
rect 22704 36700 22710 36712
rect 22741 36703 22799 36709
rect 22741 36700 22753 36703
rect 22704 36672 22753 36700
rect 22704 36660 22710 36672
rect 22741 36669 22753 36672
rect 22787 36669 22799 36703
rect 25498 36700 25504 36712
rect 22741 36663 22799 36669
rect 22848 36672 25504 36700
rect 18472 36604 18644 36632
rect 18472 36592 18478 36604
rect 20714 36592 20720 36644
rect 20772 36632 20778 36644
rect 21358 36632 21364 36644
rect 20772 36604 21364 36632
rect 20772 36592 20778 36604
rect 21358 36592 21364 36604
rect 21416 36632 21422 36644
rect 22848 36632 22876 36672
rect 25498 36660 25504 36672
rect 25556 36660 25562 36712
rect 21416 36604 22876 36632
rect 21416 36592 21422 36604
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 3418 36564 3424 36576
rect 1627 36536 3424 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 3418 36524 3424 36536
rect 3476 36524 3482 36576
rect 7190 36524 7196 36576
rect 7248 36564 7254 36576
rect 9769 36567 9827 36573
rect 9769 36564 9781 36567
rect 7248 36536 9781 36564
rect 7248 36524 7254 36536
rect 9769 36533 9781 36536
rect 9815 36533 9827 36567
rect 9769 36527 9827 36533
rect 9950 36524 9956 36576
rect 10008 36564 10014 36576
rect 11149 36567 11207 36573
rect 11149 36564 11161 36567
rect 10008 36536 11161 36564
rect 10008 36524 10014 36536
rect 11149 36533 11161 36536
rect 11195 36533 11207 36567
rect 11149 36527 11207 36533
rect 16298 36524 16304 36576
rect 16356 36564 16362 36576
rect 17037 36567 17095 36573
rect 17037 36564 17049 36567
rect 16356 36536 17049 36564
rect 16356 36524 16362 36536
rect 17037 36533 17049 36536
rect 17083 36533 17095 36567
rect 17037 36527 17095 36533
rect 20622 36524 20628 36576
rect 20680 36564 20686 36576
rect 22462 36564 22468 36576
rect 20680 36536 22468 36564
rect 20680 36524 20686 36536
rect 22462 36524 22468 36536
rect 22520 36564 22526 36576
rect 22830 36564 22836 36576
rect 22520 36536 22836 36564
rect 22520 36524 22526 36536
rect 22830 36524 22836 36536
rect 22888 36524 22894 36576
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 24489 36567 24547 36573
rect 24489 36564 24501 36567
rect 23532 36536 24501 36564
rect 23532 36524 23538 36536
rect 24489 36533 24501 36536
rect 24535 36533 24547 36567
rect 24489 36527 24547 36533
rect 24854 36524 24860 36576
rect 24912 36564 24918 36576
rect 25133 36567 25191 36573
rect 25133 36564 25145 36567
rect 24912 36536 25145 36564
rect 24912 36524 24918 36536
rect 25133 36533 25145 36536
rect 25179 36533 25191 36567
rect 25133 36527 25191 36533
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7834 36320 7840 36372
rect 7892 36320 7898 36372
rect 9030 36360 9036 36372
rect 8496 36332 9036 36360
rect 8496 36292 8524 36332
rect 9030 36320 9036 36332
rect 9088 36320 9094 36372
rect 12526 36320 12532 36372
rect 12584 36360 12590 36372
rect 13078 36360 13084 36372
rect 12584 36332 13084 36360
rect 12584 36320 12590 36332
rect 13078 36320 13084 36332
rect 13136 36320 13142 36372
rect 15933 36363 15991 36369
rect 15933 36329 15945 36363
rect 15979 36360 15991 36363
rect 18598 36360 18604 36372
rect 15979 36332 18604 36360
rect 15979 36329 15991 36332
rect 15933 36323 15991 36329
rect 18598 36320 18604 36332
rect 18656 36320 18662 36372
rect 19904 36332 20208 36360
rect 7484 36264 8524 36292
rect 6365 36227 6423 36233
rect 6365 36193 6377 36227
rect 6411 36224 6423 36227
rect 7484 36224 7512 36264
rect 8570 36252 8576 36304
rect 8628 36292 8634 36304
rect 8754 36292 8760 36304
rect 8628 36264 8760 36292
rect 8628 36252 8634 36264
rect 8754 36252 8760 36264
rect 8812 36292 8818 36304
rect 8812 36264 16436 36292
rect 8812 36252 8818 36264
rect 6411 36196 7512 36224
rect 6411 36193 6423 36196
rect 6365 36187 6423 36193
rect 7558 36184 7564 36236
rect 7616 36224 7622 36236
rect 9861 36227 9919 36233
rect 9861 36224 9873 36227
rect 7616 36196 9873 36224
rect 7616 36184 7622 36196
rect 9861 36193 9873 36196
rect 9907 36193 9919 36227
rect 9861 36187 9919 36193
rect 12710 36184 12716 36236
rect 12768 36224 12774 36236
rect 16408 36233 16436 36264
rect 16758 36252 16764 36304
rect 16816 36292 16822 36304
rect 17129 36295 17187 36301
rect 17129 36292 17141 36295
rect 16816 36264 17141 36292
rect 16816 36252 16822 36264
rect 17129 36261 17141 36264
rect 17175 36261 17187 36295
rect 18690 36292 18696 36304
rect 17129 36255 17187 36261
rect 17604 36264 18696 36292
rect 12989 36227 13047 36233
rect 12989 36224 13001 36227
rect 12768 36196 13001 36224
rect 12768 36184 12774 36196
rect 12989 36193 13001 36196
rect 13035 36193 13047 36227
rect 12989 36187 13047 36193
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36193 16451 36227
rect 16393 36187 16451 36193
rect 16577 36227 16635 36233
rect 16577 36193 16589 36227
rect 16623 36224 16635 36227
rect 17604 36224 17632 36264
rect 18690 36252 18696 36264
rect 18748 36252 18754 36304
rect 16623 36196 17632 36224
rect 16623 36193 16635 36196
rect 16577 36187 16635 36193
rect 17678 36184 17684 36236
rect 17736 36184 17742 36236
rect 4982 36116 4988 36168
rect 5040 36156 5046 36168
rect 6086 36156 6092 36168
rect 5040 36128 6092 36156
rect 5040 36116 5046 36128
rect 6086 36116 6092 36128
rect 6144 36116 6150 36168
rect 9125 36159 9183 36165
rect 9125 36125 9137 36159
rect 9171 36156 9183 36159
rect 11057 36159 11115 36165
rect 11057 36156 11069 36159
rect 9171 36128 11069 36156
rect 9171 36125 9183 36128
rect 9125 36119 9183 36125
rect 11057 36125 11069 36128
rect 11103 36156 11115 36159
rect 11422 36156 11428 36168
rect 11103 36128 11428 36156
rect 11103 36125 11115 36128
rect 11057 36119 11115 36125
rect 11422 36116 11428 36128
rect 11480 36156 11486 36168
rect 12897 36159 12955 36165
rect 11480 36128 12434 36156
rect 11480 36116 11486 36128
rect 6822 36088 6828 36100
rect 6748 36060 6828 36088
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 6748 36020 6776 36060
rect 6822 36048 6828 36060
rect 6880 36048 6886 36100
rect 11790 36048 11796 36100
rect 11848 36048 11854 36100
rect 12406 36088 12434 36128
rect 12897 36125 12909 36159
rect 12943 36156 12955 36159
rect 13354 36156 13360 36168
rect 12943 36128 13360 36156
rect 12943 36125 12955 36128
rect 12897 36119 12955 36125
rect 13354 36116 13360 36128
rect 13412 36116 13418 36168
rect 15194 36116 15200 36168
rect 15252 36156 15258 36168
rect 15381 36159 15439 36165
rect 15381 36156 15393 36159
rect 15252 36128 15393 36156
rect 15252 36116 15258 36128
rect 15381 36125 15393 36128
rect 15427 36125 15439 36159
rect 15381 36119 15439 36125
rect 16298 36116 16304 36168
rect 16356 36116 16362 36168
rect 17497 36159 17555 36165
rect 17497 36125 17509 36159
rect 17543 36156 17555 36159
rect 19904 36156 19932 36332
rect 19981 36295 20039 36301
rect 19981 36261 19993 36295
rect 20027 36261 20039 36295
rect 20180 36292 20208 36332
rect 21450 36320 21456 36372
rect 21508 36320 21514 36372
rect 21910 36320 21916 36372
rect 21968 36360 21974 36372
rect 22738 36360 22744 36372
rect 21968 36332 22744 36360
rect 21968 36320 21974 36332
rect 22738 36320 22744 36332
rect 22796 36320 22802 36372
rect 22830 36320 22836 36372
rect 22888 36360 22894 36372
rect 23750 36360 23756 36372
rect 22888 36332 23756 36360
rect 22888 36320 22894 36332
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 21266 36292 21272 36304
rect 20180 36264 21272 36292
rect 19981 36255 20039 36261
rect 17543 36128 19932 36156
rect 19996 36156 20024 36255
rect 21266 36252 21272 36264
rect 21324 36292 21330 36304
rect 25133 36295 25191 36301
rect 25133 36292 25145 36295
rect 21324 36264 25145 36292
rect 21324 36252 21330 36264
rect 25133 36261 25145 36264
rect 25179 36261 25191 36295
rect 25133 36255 25191 36261
rect 20622 36184 20628 36236
rect 20680 36184 20686 36236
rect 21726 36184 21732 36236
rect 21784 36224 21790 36236
rect 22005 36227 22063 36233
rect 22005 36224 22017 36227
rect 21784 36196 22017 36224
rect 21784 36184 21790 36196
rect 22005 36193 22017 36196
rect 22051 36224 22063 36227
rect 23474 36224 23480 36236
rect 22051 36196 23480 36224
rect 22051 36193 22063 36196
rect 22005 36187 22063 36193
rect 23474 36184 23480 36196
rect 23532 36184 23538 36236
rect 23658 36184 23664 36236
rect 23716 36224 23722 36236
rect 23753 36227 23811 36233
rect 23753 36224 23765 36227
rect 23716 36196 23765 36224
rect 23716 36184 23722 36196
rect 23753 36193 23765 36196
rect 23799 36193 23811 36227
rect 23753 36187 23811 36193
rect 23937 36227 23995 36233
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24210 36224 24216 36236
rect 23983 36196 24216 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24210 36184 24216 36196
rect 24268 36184 24274 36236
rect 25038 36156 25044 36168
rect 19996 36128 25044 36156
rect 17543 36125 17555 36128
rect 17497 36119 17555 36125
rect 25038 36116 25044 36128
rect 25096 36116 25102 36168
rect 25317 36159 25375 36165
rect 25317 36125 25329 36159
rect 25363 36156 25375 36159
rect 25498 36156 25504 36168
rect 25363 36128 25504 36156
rect 25363 36125 25375 36128
rect 25317 36119 25375 36125
rect 25498 36116 25504 36128
rect 25556 36116 25562 36168
rect 16022 36088 16028 36100
rect 12406 36060 16028 36088
rect 16022 36048 16028 36060
rect 16080 36048 16086 36100
rect 17586 36048 17592 36100
rect 17644 36048 17650 36100
rect 19058 36048 19064 36100
rect 19116 36088 19122 36100
rect 19242 36088 19248 36100
rect 19116 36060 19248 36088
rect 19116 36048 19122 36060
rect 19242 36048 19248 36060
rect 19300 36048 19306 36100
rect 20346 36048 20352 36100
rect 20404 36048 20410 36100
rect 21174 36048 21180 36100
rect 21232 36088 21238 36100
rect 21913 36091 21971 36097
rect 21913 36088 21925 36091
rect 21232 36060 21925 36088
rect 21232 36048 21238 36060
rect 21913 36057 21925 36060
rect 21959 36088 21971 36091
rect 22002 36088 22008 36100
rect 21959 36060 22008 36088
rect 21959 36057 21971 36060
rect 21913 36051 21971 36057
rect 22002 36048 22008 36060
rect 22060 36048 22066 36100
rect 22094 36048 22100 36100
rect 22152 36088 22158 36100
rect 24118 36088 24124 36100
rect 22152 36060 24124 36088
rect 22152 36048 22158 36060
rect 24118 36048 24124 36060
rect 24176 36048 24182 36100
rect 5592 35992 6776 36020
rect 5592 35980 5598 35992
rect 8294 35980 8300 36032
rect 8352 36020 8358 36032
rect 9674 36020 9680 36032
rect 8352 35992 9680 36020
rect 8352 35980 8358 35992
rect 9674 35980 9680 35992
rect 9732 35980 9738 36032
rect 12434 35980 12440 36032
rect 12492 35980 12498 36032
rect 12805 36023 12863 36029
rect 12805 35989 12817 36023
rect 12851 36020 12863 36023
rect 15286 36020 15292 36032
rect 12851 35992 15292 36020
rect 12851 35989 12863 35992
rect 12805 35983 12863 35989
rect 15286 35980 15292 35992
rect 15344 35980 15350 36032
rect 18506 35980 18512 36032
rect 18564 36020 18570 36032
rect 19334 36020 19340 36032
rect 18564 35992 19340 36020
rect 18564 35980 18570 35992
rect 19334 35980 19340 35992
rect 19392 36020 19398 36032
rect 20441 36023 20499 36029
rect 20441 36020 20453 36023
rect 19392 35992 20453 36020
rect 19392 35980 19398 35992
rect 20441 35989 20453 35992
rect 20487 36020 20499 36023
rect 20714 36020 20720 36032
rect 20487 35992 20720 36020
rect 20487 35989 20499 35992
rect 20441 35983 20499 35989
rect 20714 35980 20720 35992
rect 20772 35980 20778 36032
rect 20806 35980 20812 36032
rect 20864 36020 20870 36032
rect 21821 36023 21879 36029
rect 21821 36020 21833 36023
rect 20864 35992 21833 36020
rect 20864 35980 20870 35992
rect 21821 35989 21833 35992
rect 21867 36020 21879 36023
rect 22370 36020 22376 36032
rect 21867 35992 22376 36020
rect 21867 35989 21879 35992
rect 21821 35983 21879 35989
rect 22370 35980 22376 35992
rect 22428 35980 22434 36032
rect 22830 35980 22836 36032
rect 22888 36020 22894 36032
rect 23293 36023 23351 36029
rect 23293 36020 23305 36023
rect 22888 35992 23305 36020
rect 22888 35980 22894 35992
rect 23293 35989 23305 35992
rect 23339 35989 23351 36023
rect 23293 35983 23351 35989
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5997 35819 6055 35825
rect 5997 35785 6009 35819
rect 6043 35816 6055 35819
rect 7006 35816 7012 35828
rect 6043 35788 7012 35816
rect 6043 35785 6055 35788
rect 5997 35779 6055 35785
rect 7006 35776 7012 35788
rect 7064 35776 7070 35828
rect 9582 35776 9588 35828
rect 9640 35816 9646 35828
rect 11149 35819 11207 35825
rect 11149 35816 11161 35819
rect 9640 35788 11161 35816
rect 9640 35776 9646 35788
rect 11149 35785 11161 35788
rect 11195 35785 11207 35819
rect 11149 35779 11207 35785
rect 5534 35708 5540 35760
rect 5592 35708 5598 35760
rect 9674 35708 9680 35760
rect 9732 35748 9738 35760
rect 10134 35748 10140 35760
rect 9732 35720 10140 35748
rect 9732 35708 9738 35720
rect 10134 35708 10140 35720
rect 10192 35708 10198 35760
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35581 4307 35615
rect 4249 35575 4307 35581
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 6822 35612 6828 35624
rect 4571 35584 6828 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 4264 35476 4292 35575
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 9214 35572 9220 35624
rect 9272 35612 9278 35624
rect 9401 35615 9459 35621
rect 9401 35612 9413 35615
rect 9272 35584 9413 35612
rect 9272 35572 9278 35584
rect 9401 35581 9413 35584
rect 9447 35581 9459 35615
rect 9401 35575 9459 35581
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 10686 35612 10692 35624
rect 9723 35584 10692 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 10686 35572 10692 35584
rect 10744 35612 10750 35624
rect 11054 35612 11060 35624
rect 10744 35584 11060 35612
rect 10744 35572 10750 35584
rect 11054 35572 11060 35584
rect 11112 35572 11118 35624
rect 4982 35476 4988 35488
rect 4212 35448 4988 35476
rect 4212 35436 4218 35448
rect 4982 35436 4988 35448
rect 5040 35436 5046 35488
rect 11164 35476 11192 35779
rect 12802 35776 12808 35828
rect 12860 35816 12866 35828
rect 13541 35819 13599 35825
rect 13541 35816 13553 35819
rect 12860 35788 13553 35816
rect 12860 35776 12866 35788
rect 13541 35785 13553 35788
rect 13587 35785 13599 35819
rect 13541 35779 13599 35785
rect 13630 35776 13636 35828
rect 13688 35816 13694 35828
rect 14461 35819 14519 35825
rect 14461 35816 14473 35819
rect 13688 35788 14473 35816
rect 13688 35776 13694 35788
rect 14461 35785 14473 35788
rect 14507 35785 14519 35819
rect 14461 35779 14519 35785
rect 15102 35776 15108 35828
rect 15160 35816 15166 35828
rect 15197 35819 15255 35825
rect 15197 35816 15209 35819
rect 15160 35788 15209 35816
rect 15160 35776 15166 35788
rect 15197 35785 15209 35788
rect 15243 35785 15255 35819
rect 15197 35779 15255 35785
rect 16850 35776 16856 35828
rect 16908 35776 16914 35828
rect 18598 35816 18604 35828
rect 16960 35788 18604 35816
rect 14369 35751 14427 35757
rect 14369 35717 14381 35751
rect 14415 35748 14427 35751
rect 16960 35748 16988 35788
rect 18598 35776 18604 35788
rect 18656 35776 18662 35828
rect 20162 35816 20168 35828
rect 18708 35788 20168 35816
rect 14415 35720 16988 35748
rect 14415 35717 14427 35720
rect 14369 35711 14427 35717
rect 17034 35708 17040 35760
rect 17092 35748 17098 35760
rect 18708 35748 18736 35788
rect 20162 35776 20168 35788
rect 20220 35776 20226 35828
rect 17092 35720 18736 35748
rect 17092 35708 17098 35720
rect 13354 35680 13360 35692
rect 13202 35652 13360 35680
rect 13354 35640 13360 35652
rect 13412 35640 13418 35692
rect 15565 35683 15623 35689
rect 15565 35680 15577 35683
rect 14568 35652 15577 35680
rect 11790 35572 11796 35624
rect 11848 35572 11854 35624
rect 12069 35615 12127 35621
rect 12069 35581 12081 35615
rect 12115 35612 12127 35615
rect 14182 35612 14188 35624
rect 12115 35584 14188 35612
rect 12115 35581 12127 35584
rect 12069 35575 12127 35581
rect 14182 35572 14188 35584
rect 14240 35572 14246 35624
rect 13078 35504 13084 35556
rect 13136 35544 13142 35556
rect 14568 35544 14596 35652
rect 15565 35649 15577 35652
rect 15611 35680 15623 35683
rect 16298 35680 16304 35692
rect 15611 35652 16304 35680
rect 15611 35649 15623 35652
rect 15565 35643 15623 35649
rect 16298 35640 16304 35652
rect 16356 35640 16362 35692
rect 18616 35689 18644 35720
rect 18782 35708 18788 35760
rect 18840 35748 18846 35760
rect 18877 35751 18935 35757
rect 18877 35748 18889 35751
rect 18840 35720 18889 35748
rect 18840 35708 18846 35720
rect 18877 35717 18889 35720
rect 18923 35717 18935 35751
rect 18877 35711 18935 35717
rect 19334 35708 19340 35760
rect 19392 35708 19398 35760
rect 23474 35708 23480 35760
rect 23532 35708 23538 35760
rect 24486 35708 24492 35760
rect 24544 35708 24550 35760
rect 17221 35683 17279 35689
rect 17221 35649 17233 35683
rect 17267 35680 17279 35683
rect 18601 35683 18659 35689
rect 17267 35652 18552 35680
rect 17267 35649 17279 35652
rect 17221 35643 17279 35649
rect 14645 35615 14703 35621
rect 14645 35581 14657 35615
rect 14691 35612 14703 35615
rect 15286 35612 15292 35624
rect 14691 35584 15292 35612
rect 14691 35581 14703 35584
rect 14645 35575 14703 35581
rect 15286 35572 15292 35584
rect 15344 35572 15350 35624
rect 15657 35615 15715 35621
rect 15657 35581 15669 35615
rect 15703 35581 15715 35615
rect 15657 35575 15715 35581
rect 15841 35615 15899 35621
rect 15841 35581 15853 35615
rect 15887 35612 15899 35615
rect 16390 35612 16396 35624
rect 15887 35584 16396 35612
rect 15887 35581 15899 35584
rect 15841 35575 15899 35581
rect 13136 35516 14596 35544
rect 15672 35544 15700 35575
rect 16390 35572 16396 35584
rect 16448 35572 16454 35624
rect 17310 35572 17316 35624
rect 17368 35572 17374 35624
rect 17405 35615 17463 35621
rect 17405 35581 17417 35615
rect 17451 35581 17463 35615
rect 18524 35612 18552 35652
rect 18601 35649 18613 35683
rect 18647 35649 18659 35683
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 18601 35643 18659 35649
rect 20640 35652 22048 35680
rect 18524 35584 18736 35612
rect 17405 35575 17463 35581
rect 17126 35544 17132 35556
rect 15672 35516 17132 35544
rect 13136 35504 13142 35516
rect 17126 35504 17132 35516
rect 17184 35504 17190 35556
rect 13446 35476 13452 35488
rect 11164 35448 13452 35476
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 13998 35436 14004 35488
rect 14056 35436 14062 35488
rect 14642 35436 14648 35488
rect 14700 35476 14706 35488
rect 17420 35476 17448 35575
rect 14700 35448 17448 35476
rect 18708 35476 18736 35584
rect 19242 35572 19248 35624
rect 19300 35612 19306 35624
rect 20640 35612 20668 35652
rect 19300 35584 20668 35612
rect 19300 35572 19306 35584
rect 22020 35544 22048 35652
rect 22204 35652 22385 35680
rect 22204 35544 22232 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 22465 35683 22523 35689
rect 22465 35649 22477 35683
rect 22511 35680 22523 35683
rect 22738 35680 22744 35692
rect 22511 35652 22744 35680
rect 22511 35649 22523 35652
rect 22465 35643 22523 35649
rect 22738 35640 22744 35652
rect 22796 35640 22802 35692
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 22646 35572 22652 35624
rect 22704 35612 22710 35624
rect 23201 35615 23259 35621
rect 23201 35612 23213 35615
rect 22704 35584 23213 35612
rect 22704 35572 22710 35584
rect 23201 35581 23213 35584
rect 23247 35581 23259 35615
rect 23201 35575 23259 35581
rect 22020 35516 22232 35544
rect 19334 35476 19340 35488
rect 18708 35448 19340 35476
rect 14700 35436 14706 35448
rect 19334 35436 19340 35448
rect 19392 35436 19398 35488
rect 20349 35479 20407 35485
rect 20349 35445 20361 35479
rect 20395 35476 20407 35479
rect 21082 35476 21088 35488
rect 20395 35448 21088 35476
rect 20395 35445 20407 35448
rect 20349 35439 20407 35445
rect 21082 35436 21088 35448
rect 21140 35436 21146 35488
rect 22005 35479 22063 35485
rect 22005 35445 22017 35479
rect 22051 35476 22063 35479
rect 22738 35476 22744 35488
rect 22051 35448 22744 35476
rect 22051 35445 22063 35448
rect 22005 35439 22063 35445
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 23290 35436 23296 35488
rect 23348 35476 23354 35488
rect 24949 35479 25007 35485
rect 24949 35476 24961 35479
rect 23348 35448 24961 35476
rect 23348 35436 23354 35448
rect 24949 35445 24961 35448
rect 24995 35445 25007 35479
rect 24949 35439 25007 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 7098 35232 7104 35284
rect 7156 35272 7162 35284
rect 7653 35275 7711 35281
rect 7653 35272 7665 35275
rect 7156 35244 7665 35272
rect 7156 35232 7162 35244
rect 7653 35241 7665 35244
rect 7699 35241 7711 35275
rect 7653 35235 7711 35241
rect 9585 35275 9643 35281
rect 9585 35241 9597 35275
rect 9631 35272 9643 35275
rect 10042 35272 10048 35284
rect 9631 35244 10048 35272
rect 9631 35241 9643 35244
rect 9585 35235 9643 35241
rect 10042 35232 10048 35244
rect 10100 35232 10106 35284
rect 14829 35275 14887 35281
rect 14829 35241 14841 35275
rect 14875 35272 14887 35275
rect 15562 35272 15568 35284
rect 14875 35244 15568 35272
rect 14875 35241 14887 35244
rect 14829 35235 14887 35241
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 17310 35232 17316 35284
rect 17368 35272 17374 35284
rect 19702 35272 19708 35284
rect 17368 35244 19708 35272
rect 17368 35232 17374 35244
rect 19702 35232 19708 35244
rect 19760 35272 19766 35284
rect 21542 35272 21548 35284
rect 19760 35244 21548 35272
rect 19760 35232 19766 35244
rect 21542 35232 21548 35244
rect 21600 35232 21606 35284
rect 22833 35275 22891 35281
rect 22833 35241 22845 35275
rect 22879 35272 22891 35275
rect 23658 35272 23664 35284
rect 22879 35244 23664 35272
rect 22879 35241 22891 35244
rect 22833 35235 22891 35241
rect 23658 35232 23664 35244
rect 23716 35232 23722 35284
rect 7282 35204 7288 35216
rect 6840 35176 7288 35204
rect 5537 35139 5595 35145
rect 5537 35105 5549 35139
rect 5583 35136 5595 35139
rect 6840 35136 6868 35176
rect 7282 35164 7288 35176
rect 7340 35204 7346 35216
rect 7558 35204 7564 35216
rect 7340 35176 7564 35204
rect 7340 35164 7346 35176
rect 7558 35164 7564 35176
rect 7616 35164 7622 35216
rect 9214 35164 9220 35216
rect 9272 35204 9278 35216
rect 11790 35204 11796 35216
rect 9272 35176 11796 35204
rect 9272 35164 9278 35176
rect 11790 35164 11796 35176
rect 11848 35204 11854 35216
rect 11848 35176 12020 35204
rect 11848 35164 11854 35176
rect 5583 35108 6868 35136
rect 5583 35105 5595 35108
rect 5537 35099 5595 35105
rect 6914 35096 6920 35148
rect 6972 35136 6978 35148
rect 8205 35139 8263 35145
rect 8205 35136 8217 35139
rect 6972 35108 8217 35136
rect 6972 35096 6978 35108
rect 8205 35105 8217 35108
rect 8251 35105 8263 35139
rect 8205 35099 8263 35105
rect 9582 35096 9588 35148
rect 9640 35136 9646 35148
rect 10137 35139 10195 35145
rect 10137 35136 10149 35139
rect 9640 35108 10149 35136
rect 9640 35096 9646 35108
rect 10137 35105 10149 35108
rect 10183 35105 10195 35139
rect 10137 35099 10195 35105
rect 4982 35028 4988 35080
rect 5040 35068 5046 35080
rect 5261 35071 5319 35077
rect 5261 35068 5273 35071
rect 5040 35040 5273 35068
rect 5040 35028 5046 35040
rect 5261 35037 5273 35040
rect 5307 35037 5319 35071
rect 5261 35031 5319 35037
rect 9950 35028 9956 35080
rect 10008 35028 10014 35080
rect 11992 35077 12020 35176
rect 13446 35164 13452 35216
rect 13504 35204 13510 35216
rect 13504 35176 16712 35204
rect 13504 35164 13510 35176
rect 12253 35139 12311 35145
rect 12253 35105 12265 35139
rect 12299 35136 12311 35139
rect 12299 35108 13584 35136
rect 12299 35105 12311 35108
rect 12253 35099 12311 35105
rect 11977 35071 12035 35077
rect 11977 35037 11989 35071
rect 12023 35037 12035 35071
rect 11977 35031 12035 35037
rect 13354 35028 13360 35080
rect 13412 35028 13418 35080
rect 13556 35068 13584 35108
rect 13630 35096 13636 35148
rect 13688 35136 13694 35148
rect 15289 35139 15347 35145
rect 15289 35136 15301 35139
rect 13688 35108 15301 35136
rect 13688 35096 13694 35108
rect 15289 35105 15301 35108
rect 15335 35105 15347 35139
rect 15289 35099 15347 35105
rect 15473 35139 15531 35145
rect 15473 35105 15485 35139
rect 15519 35136 15531 35139
rect 16574 35136 16580 35148
rect 15519 35108 16580 35136
rect 15519 35105 15531 35108
rect 15473 35099 15531 35105
rect 16574 35096 16580 35108
rect 16632 35096 16638 35148
rect 16684 35136 16712 35176
rect 17126 35164 17132 35216
rect 17184 35204 17190 35216
rect 17954 35204 17960 35216
rect 17184 35176 17960 35204
rect 17184 35164 17190 35176
rect 17954 35164 17960 35176
rect 18012 35164 18018 35216
rect 18141 35207 18199 35213
rect 18141 35173 18153 35207
rect 18187 35204 18199 35207
rect 18966 35204 18972 35216
rect 18187 35176 18972 35204
rect 18187 35173 18199 35176
rect 18141 35167 18199 35173
rect 18966 35164 18972 35176
rect 19024 35164 19030 35216
rect 19334 35164 19340 35216
rect 19392 35204 19398 35216
rect 25133 35207 25191 35213
rect 25133 35204 25145 35207
rect 19392 35176 25145 35204
rect 19392 35164 19398 35176
rect 25133 35173 25145 35176
rect 25179 35173 25191 35207
rect 25133 35167 25191 35173
rect 18693 35139 18751 35145
rect 18693 35136 18705 35139
rect 16684 35108 18705 35136
rect 18693 35105 18705 35108
rect 18739 35105 18751 35139
rect 18693 35099 18751 35105
rect 19610 35096 19616 35148
rect 19668 35136 19674 35148
rect 20533 35139 20591 35145
rect 20533 35136 20545 35139
rect 19668 35108 20545 35136
rect 19668 35096 19674 35108
rect 20533 35105 20545 35108
rect 20579 35105 20591 35139
rect 20533 35099 20591 35105
rect 20714 35096 20720 35148
rect 20772 35136 20778 35148
rect 22094 35136 22100 35148
rect 20772 35108 22100 35136
rect 20772 35096 20778 35108
rect 22094 35096 22100 35108
rect 22152 35096 22158 35148
rect 22462 35096 22468 35148
rect 22520 35136 22526 35148
rect 23198 35136 23204 35148
rect 22520 35108 23204 35136
rect 22520 35096 22526 35108
rect 23198 35096 23204 35108
rect 23256 35096 23262 35148
rect 23290 35096 23296 35148
rect 23348 35136 23354 35148
rect 23385 35139 23443 35145
rect 23385 35136 23397 35139
rect 23348 35108 23397 35136
rect 23348 35096 23354 35108
rect 23385 35105 23397 35108
rect 23431 35105 23443 35139
rect 23385 35099 23443 35105
rect 13814 35068 13820 35080
rect 13556 35040 13820 35068
rect 13814 35028 13820 35040
rect 13872 35068 13878 35080
rect 14826 35068 14832 35080
rect 13872 35040 14832 35068
rect 13872 35028 13878 35040
rect 14826 35028 14832 35040
rect 14884 35028 14890 35080
rect 15194 35028 15200 35080
rect 15252 35028 15258 35080
rect 18601 35071 18659 35077
rect 18601 35037 18613 35071
rect 18647 35068 18659 35071
rect 20349 35071 20407 35077
rect 20349 35068 20361 35071
rect 18647 35040 20361 35068
rect 18647 35037 18659 35040
rect 18601 35031 18659 35037
rect 20349 35037 20361 35040
rect 20395 35068 20407 35071
rect 25130 35068 25136 35080
rect 20395 35040 25136 35068
rect 20395 35037 20407 35040
rect 20349 35031 20407 35037
rect 25130 35028 25136 35040
rect 25188 35028 25194 35080
rect 25317 35071 25375 35077
rect 25317 35037 25329 35071
rect 25363 35068 25375 35071
rect 25406 35068 25412 35080
rect 25363 35040 25412 35068
rect 25363 35037 25375 35040
rect 25317 35031 25375 35037
rect 25406 35028 25412 35040
rect 25464 35028 25470 35080
rect 5534 34960 5540 35012
rect 5592 35000 5598 35012
rect 5592 34972 6026 35000
rect 5592 34960 5598 34972
rect 6822 34960 6828 35012
rect 6880 35000 6886 35012
rect 10318 35000 10324 35012
rect 6880 34972 10324 35000
rect 6880 34960 6886 34972
rect 7024 34941 7052 34972
rect 10318 34960 10324 34972
rect 10376 34960 10382 35012
rect 7009 34935 7067 34941
rect 7009 34901 7021 34935
rect 7055 34901 7067 34935
rect 7009 34895 7067 34901
rect 7834 34892 7840 34944
rect 7892 34932 7898 34944
rect 8021 34935 8079 34941
rect 8021 34932 8033 34935
rect 7892 34904 8033 34932
rect 7892 34892 7898 34904
rect 8021 34901 8033 34904
rect 8067 34901 8079 34935
rect 8021 34895 8079 34901
rect 8113 34935 8171 34941
rect 8113 34901 8125 34935
rect 8159 34932 8171 34935
rect 9582 34932 9588 34944
rect 8159 34904 9588 34932
rect 8159 34901 8171 34904
rect 8113 34895 8171 34901
rect 9582 34892 9588 34904
rect 9640 34892 9646 34944
rect 10042 34892 10048 34944
rect 10100 34892 10106 34944
rect 10134 34892 10140 34944
rect 10192 34932 10198 34944
rect 13372 34932 13400 35028
rect 18690 34960 18696 35012
rect 18748 35000 18754 35012
rect 18748 34972 20024 35000
rect 18748 34960 18754 34972
rect 10192 34904 13400 34932
rect 13725 34935 13783 34941
rect 10192 34892 10198 34904
rect 13725 34901 13737 34935
rect 13771 34932 13783 34935
rect 14182 34932 14188 34944
rect 13771 34904 14188 34932
rect 13771 34901 13783 34904
rect 13725 34895 13783 34901
rect 14182 34892 14188 34904
rect 14240 34892 14246 34944
rect 18509 34935 18567 34941
rect 18509 34901 18521 34935
rect 18555 34932 18567 34935
rect 18874 34932 18880 34944
rect 18555 34904 18880 34932
rect 18555 34901 18567 34904
rect 18509 34895 18567 34901
rect 18874 34892 18880 34904
rect 18932 34892 18938 34944
rect 19996 34941 20024 34972
rect 20070 34960 20076 35012
rect 20128 35000 20134 35012
rect 20441 35003 20499 35009
rect 20441 35000 20453 35003
rect 20128 34972 20453 35000
rect 20128 34960 20134 34972
rect 20441 34969 20453 34972
rect 20487 34969 20499 35003
rect 20441 34963 20499 34969
rect 20714 34960 20720 35012
rect 20772 35000 20778 35012
rect 23293 35003 23351 35009
rect 23293 35000 23305 35003
rect 20772 34972 23305 35000
rect 20772 34960 20778 34972
rect 23293 34969 23305 34972
rect 23339 34969 23351 35003
rect 23293 34963 23351 34969
rect 19981 34935 20039 34941
rect 19981 34901 19993 34935
rect 20027 34901 20039 34935
rect 19981 34895 20039 34901
rect 23198 34892 23204 34944
rect 23256 34892 23262 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 3326 34728 3332 34740
rect 1627 34700 3332 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 3326 34688 3332 34700
rect 3384 34688 3390 34740
rect 4154 34688 4160 34740
rect 4212 34688 4218 34740
rect 5258 34688 5264 34740
rect 5316 34688 5322 34740
rect 6546 34728 6552 34740
rect 5552 34700 6552 34728
rect 4172 34660 4200 34688
rect 5552 34672 5580 34700
rect 6546 34688 6552 34700
rect 6604 34728 6610 34740
rect 6604 34700 7420 34728
rect 6604 34688 6610 34700
rect 5534 34660 5540 34672
rect 3528 34632 4200 34660
rect 5014 34632 5540 34660
rect 1762 34552 1768 34604
rect 1820 34552 1826 34604
rect 3528 34601 3556 34632
rect 5534 34620 5540 34632
rect 5592 34620 5598 34672
rect 7006 34620 7012 34672
rect 7064 34620 7070 34672
rect 7392 34660 7420 34700
rect 7650 34688 7656 34740
rect 7708 34728 7714 34740
rect 9033 34731 9091 34737
rect 9033 34728 9045 34731
rect 7708 34700 9045 34728
rect 7708 34688 7714 34700
rect 9033 34697 9045 34700
rect 9079 34697 9091 34731
rect 9033 34691 9091 34697
rect 9493 34731 9551 34737
rect 9493 34697 9505 34731
rect 9539 34728 9551 34731
rect 11974 34728 11980 34740
rect 9539 34700 11980 34728
rect 9539 34697 9551 34700
rect 9493 34691 9551 34697
rect 11974 34688 11980 34700
rect 12032 34688 12038 34740
rect 12066 34688 12072 34740
rect 12124 34728 12130 34740
rect 14093 34731 14151 34737
rect 14093 34728 14105 34731
rect 12124 34700 14105 34728
rect 12124 34688 12130 34700
rect 14093 34697 14105 34700
rect 14139 34697 14151 34731
rect 14093 34691 14151 34697
rect 14461 34731 14519 34737
rect 14461 34697 14473 34731
rect 14507 34728 14519 34731
rect 14507 34700 19564 34728
rect 14507 34697 14519 34700
rect 14461 34691 14519 34697
rect 13354 34660 13360 34672
rect 7392 34632 7498 34660
rect 13202 34632 13360 34660
rect 13354 34620 13360 34632
rect 13412 34620 13418 34672
rect 14553 34663 14611 34669
rect 14553 34629 14565 34663
rect 14599 34660 14611 34663
rect 15010 34660 15016 34672
rect 14599 34632 15016 34660
rect 14599 34629 14611 34632
rect 14553 34623 14611 34629
rect 15010 34620 15016 34632
rect 15068 34620 15074 34672
rect 17034 34660 17040 34672
rect 16868 34632 17040 34660
rect 16868 34604 16896 34632
rect 17034 34620 17040 34632
rect 17092 34620 17098 34672
rect 19058 34660 19064 34672
rect 18354 34632 19064 34660
rect 19058 34620 19064 34632
rect 19116 34620 19122 34672
rect 3513 34595 3571 34601
rect 3513 34561 3525 34595
rect 3559 34561 3571 34595
rect 3513 34555 3571 34561
rect 9401 34595 9459 34601
rect 9401 34561 9413 34595
rect 9447 34561 9459 34595
rect 9401 34555 9459 34561
rect 6733 34527 6791 34533
rect 6733 34493 6745 34527
rect 6779 34524 6791 34527
rect 6779 34496 6868 34524
rect 6779 34493 6791 34496
rect 6733 34487 6791 34493
rect 3776 34391 3834 34397
rect 3776 34357 3788 34391
rect 3822 34388 3834 34391
rect 4154 34388 4160 34400
rect 3822 34360 4160 34388
rect 3822 34357 3834 34360
rect 3776 34351 3834 34357
rect 4154 34348 4160 34360
rect 4212 34348 4218 34400
rect 6840 34388 6868 34496
rect 7650 34484 7656 34536
rect 7708 34524 7714 34536
rect 9416 34524 9444 34555
rect 11698 34552 11704 34604
rect 11756 34552 11762 34604
rect 16850 34552 16856 34604
rect 16908 34552 16914 34604
rect 19429 34595 19487 34601
rect 19429 34561 19441 34595
rect 19475 34561 19487 34595
rect 19536 34592 19564 34700
rect 21174 34688 21180 34740
rect 21232 34728 21238 34740
rect 22005 34731 22063 34737
rect 22005 34728 22017 34731
rect 21232 34700 22017 34728
rect 21232 34688 21238 34700
rect 22005 34697 22017 34700
rect 22051 34697 22063 34731
rect 22005 34691 22063 34697
rect 22373 34731 22431 34737
rect 22373 34697 22385 34731
rect 22419 34728 22431 34731
rect 23382 34728 23388 34740
rect 22419 34700 23388 34728
rect 22419 34697 22431 34700
rect 22373 34691 22431 34697
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 25038 34688 25044 34740
rect 25096 34728 25102 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 25096 34700 25145 34728
rect 25096 34688 25102 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 20990 34620 20996 34672
rect 21048 34660 21054 34672
rect 22465 34663 22523 34669
rect 22465 34660 22477 34663
rect 21048 34632 22477 34660
rect 21048 34620 21054 34632
rect 22465 34629 22477 34632
rect 22511 34629 22523 34663
rect 22465 34623 22523 34629
rect 22554 34620 22560 34672
rect 22612 34660 22618 34672
rect 24302 34660 24308 34672
rect 22612 34632 24308 34660
rect 22612 34620 22618 34632
rect 22756 34592 22784 34632
rect 24302 34620 24308 34632
rect 24360 34620 24366 34672
rect 19536 34564 22784 34592
rect 19429 34555 19487 34561
rect 7708 34496 9444 34524
rect 9585 34527 9643 34533
rect 7708 34484 7714 34496
rect 9585 34493 9597 34527
rect 9631 34493 9643 34527
rect 9585 34487 9643 34493
rect 11977 34527 12035 34533
rect 11977 34493 11989 34527
rect 12023 34524 12035 34527
rect 12618 34524 12624 34536
rect 12023 34496 12624 34524
rect 12023 34493 12035 34496
rect 11977 34487 12035 34493
rect 8294 34416 8300 34468
rect 8352 34456 8358 34468
rect 9600 34456 9628 34487
rect 12618 34484 12624 34496
rect 12676 34484 12682 34536
rect 13354 34484 13360 34536
rect 13412 34524 13418 34536
rect 13449 34527 13507 34533
rect 13449 34524 13461 34527
rect 13412 34496 13461 34524
rect 13412 34484 13418 34496
rect 13449 34493 13461 34496
rect 13495 34493 13507 34527
rect 13449 34487 13507 34493
rect 14737 34527 14795 34533
rect 14737 34493 14749 34527
rect 14783 34493 14795 34527
rect 14737 34487 14795 34493
rect 8352 34428 9628 34456
rect 14752 34456 14780 34487
rect 17126 34484 17132 34536
rect 17184 34484 17190 34536
rect 18322 34484 18328 34536
rect 18380 34524 18386 34536
rect 18601 34527 18659 34533
rect 18601 34524 18613 34527
rect 18380 34496 18613 34524
rect 18380 34484 18386 34496
rect 18601 34493 18613 34496
rect 18647 34493 18659 34527
rect 19242 34524 19248 34536
rect 18601 34487 18659 34493
rect 19076 34496 19248 34524
rect 14826 34456 14832 34468
rect 14752 34428 14832 34456
rect 8352 34416 8358 34428
rect 14826 34416 14832 34428
rect 14884 34416 14890 34468
rect 19076 34465 19104 34496
rect 19242 34484 19248 34496
rect 19300 34484 19306 34536
rect 19061 34459 19119 34465
rect 19061 34425 19073 34459
rect 19107 34425 19119 34459
rect 19061 34419 19119 34425
rect 7742 34388 7748 34400
rect 6840 34360 7748 34388
rect 7742 34348 7748 34360
rect 7800 34348 7806 34400
rect 8478 34348 8484 34400
rect 8536 34348 8542 34400
rect 14550 34348 14556 34400
rect 14608 34388 14614 34400
rect 15102 34388 15108 34400
rect 14608 34360 15108 34388
rect 14608 34348 14614 34360
rect 15102 34348 15108 34360
rect 15160 34348 15166 34400
rect 19444 34388 19472 34555
rect 23198 34552 23204 34604
rect 23256 34592 23262 34604
rect 23385 34595 23443 34601
rect 23385 34592 23397 34595
rect 23256 34564 23397 34592
rect 23256 34552 23262 34564
rect 23385 34561 23397 34564
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 19518 34484 19524 34536
rect 19576 34484 19582 34536
rect 19705 34527 19763 34533
rect 19705 34493 19717 34527
rect 19751 34524 19763 34527
rect 22557 34527 22615 34533
rect 19751 34496 20576 34524
rect 19751 34493 19763 34496
rect 19705 34487 19763 34493
rect 20441 34459 20499 34465
rect 20441 34425 20453 34459
rect 20487 34425 20499 34459
rect 20548 34456 20576 34496
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 22557 34487 22615 34493
rect 21634 34456 21640 34468
rect 20548 34428 21640 34456
rect 20441 34419 20499 34425
rect 20456 34388 20484 34419
rect 21634 34416 21640 34428
rect 21692 34416 21698 34468
rect 22462 34416 22468 34468
rect 22520 34456 22526 34468
rect 22572 34456 22600 34487
rect 22520 34428 22600 34456
rect 22520 34416 22526 34428
rect 19444 34360 20484 34388
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 4154 34144 4160 34196
rect 4212 34184 4218 34196
rect 5350 34184 5356 34196
rect 4212 34156 5356 34184
rect 4212 34144 4218 34156
rect 5350 34144 5356 34156
rect 5408 34184 5414 34196
rect 5408 34156 6684 34184
rect 5408 34144 5414 34156
rect 6656 34125 6684 34156
rect 6730 34144 6736 34196
rect 6788 34184 6794 34196
rect 6788 34156 9076 34184
rect 6788 34144 6794 34156
rect 6641 34119 6699 34125
rect 6641 34085 6653 34119
rect 6687 34116 6699 34119
rect 9048 34116 9076 34156
rect 9122 34144 9128 34196
rect 9180 34144 9186 34196
rect 11885 34187 11943 34193
rect 11885 34153 11897 34187
rect 11931 34184 11943 34187
rect 12250 34184 12256 34196
rect 11931 34156 12256 34184
rect 11931 34153 11943 34156
rect 11885 34147 11943 34153
rect 12250 34144 12256 34156
rect 12308 34144 12314 34196
rect 17126 34144 17132 34196
rect 17184 34184 17190 34196
rect 20990 34184 20996 34196
rect 17184 34156 20996 34184
rect 17184 34144 17190 34156
rect 20990 34144 20996 34156
rect 21048 34144 21054 34196
rect 11698 34116 11704 34128
rect 6687 34088 6960 34116
rect 9048 34088 11704 34116
rect 6687 34085 6699 34088
rect 6641 34079 6699 34085
rect 5169 34051 5227 34057
rect 5169 34017 5181 34051
rect 5215 34048 5227 34051
rect 6822 34048 6828 34060
rect 5215 34020 6828 34048
rect 5215 34017 5227 34020
rect 5169 34011 5227 34017
rect 6822 34008 6828 34020
rect 6880 34008 6886 34060
rect 6932 34048 6960 34088
rect 11698 34076 11704 34088
rect 11756 34116 11762 34128
rect 11756 34088 12296 34116
rect 11756 34076 11762 34088
rect 12268 34060 12296 34088
rect 12342 34076 12348 34128
rect 12400 34116 12406 34128
rect 12400 34076 12434 34116
rect 14734 34076 14740 34128
rect 14792 34116 14798 34128
rect 19886 34116 19892 34128
rect 14792 34088 19892 34116
rect 14792 34076 14798 34088
rect 19886 34076 19892 34088
rect 19944 34076 19950 34128
rect 23290 34076 23296 34128
rect 23348 34116 23354 34128
rect 24854 34116 24860 34128
rect 23348 34088 24860 34116
rect 23348 34076 23354 34088
rect 24854 34076 24860 34088
rect 24912 34076 24918 34128
rect 9677 34051 9735 34057
rect 9677 34048 9689 34051
rect 6932 34020 9689 34048
rect 9677 34017 9689 34020
rect 9723 34017 9735 34051
rect 9677 34011 9735 34017
rect 12250 34008 12256 34060
rect 12308 34008 12314 34060
rect 12406 34048 12434 34076
rect 12406 34020 12480 34048
rect 4890 33940 4896 33992
rect 4948 33940 4954 33992
rect 9585 33983 9643 33989
rect 9585 33949 9597 33983
rect 9631 33980 9643 33983
rect 12342 33980 12348 33992
rect 9631 33952 12348 33980
rect 9631 33949 9643 33952
rect 9585 33943 9643 33949
rect 12342 33940 12348 33952
rect 12400 33940 12406 33992
rect 12452 33980 12480 34020
rect 12526 34008 12532 34060
rect 12584 34048 12590 34060
rect 13446 34048 13452 34060
rect 12584 34020 13452 34048
rect 12584 34008 12590 34020
rect 13446 34008 13452 34020
rect 13504 34008 13510 34060
rect 18414 34008 18420 34060
rect 18472 34048 18478 34060
rect 19981 34051 20039 34057
rect 19981 34048 19993 34051
rect 18472 34020 19993 34048
rect 18472 34008 18478 34020
rect 19981 34017 19993 34020
rect 20027 34017 20039 34051
rect 19981 34011 20039 34017
rect 20530 34008 20536 34060
rect 20588 34048 20594 34060
rect 20993 34051 21051 34057
rect 20993 34048 21005 34051
rect 20588 34020 21005 34048
rect 20588 34008 20594 34020
rect 20993 34017 21005 34020
rect 21039 34017 21051 34051
rect 20993 34011 21051 34017
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 23624 34020 24808 34048
rect 23624 34008 23630 34020
rect 17034 33980 17040 33992
rect 12452 33952 17040 33980
rect 17034 33940 17040 33952
rect 17092 33940 17098 33992
rect 17954 33940 17960 33992
rect 18012 33980 18018 33992
rect 19797 33983 19855 33989
rect 19797 33980 19809 33983
rect 18012 33952 19809 33980
rect 18012 33940 18018 33952
rect 19797 33949 19809 33952
rect 19843 33949 19855 33983
rect 19797 33943 19855 33949
rect 5626 33872 5632 33924
rect 5684 33872 5690 33924
rect 11882 33872 11888 33924
rect 11940 33912 11946 33924
rect 11940 33884 12388 33912
rect 11940 33872 11946 33884
rect 9493 33847 9551 33853
rect 9493 33813 9505 33847
rect 9539 33844 9551 33847
rect 11974 33844 11980 33856
rect 9539 33816 11980 33844
rect 9539 33813 9551 33816
rect 9493 33807 9551 33813
rect 11974 33804 11980 33816
rect 12032 33804 12038 33856
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 12360 33853 12388 33884
rect 13262 33872 13268 33924
rect 13320 33912 13326 33924
rect 18966 33912 18972 33924
rect 13320 33884 18972 33912
rect 13320 33872 13326 33884
rect 18966 33872 18972 33884
rect 19024 33872 19030 33924
rect 19812 33912 19840 33943
rect 20346 33940 20352 33992
rect 20404 33980 20410 33992
rect 20717 33983 20775 33989
rect 20717 33980 20729 33983
rect 20404 33952 20729 33980
rect 20404 33940 20410 33952
rect 20717 33949 20729 33952
rect 20763 33949 20775 33983
rect 20717 33943 20775 33949
rect 23842 33940 23848 33992
rect 23900 33940 23906 33992
rect 24780 33989 24808 34020
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 24486 33912 24492 33924
rect 19812 33884 20852 33912
rect 22218 33884 24492 33912
rect 20824 33856 20852 33884
rect 12345 33847 12403 33853
rect 12345 33813 12357 33847
rect 12391 33813 12403 33847
rect 12345 33807 12403 33813
rect 12802 33804 12808 33856
rect 12860 33844 12866 33856
rect 13998 33844 14004 33856
rect 12860 33816 14004 33844
rect 12860 33804 12866 33816
rect 13998 33804 14004 33816
rect 14056 33804 14062 33856
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 19429 33847 19487 33853
rect 19429 33844 19441 33847
rect 16632 33816 19441 33844
rect 16632 33804 16638 33816
rect 19429 33813 19441 33816
rect 19475 33813 19487 33847
rect 19429 33807 19487 33813
rect 19794 33804 19800 33856
rect 19852 33844 19858 33856
rect 19889 33847 19947 33853
rect 19889 33844 19901 33847
rect 19852 33816 19901 33844
rect 19852 33804 19858 33816
rect 19889 33813 19901 33816
rect 19935 33813 19947 33847
rect 19889 33807 19947 33813
rect 20806 33804 20812 33856
rect 20864 33804 20870 33856
rect 21910 33804 21916 33856
rect 21968 33844 21974 33856
rect 22296 33844 22324 33884
rect 24486 33872 24492 33884
rect 24544 33872 24550 33924
rect 21968 33816 22324 33844
rect 21968 33804 21974 33816
rect 22462 33804 22468 33856
rect 22520 33804 22526 33856
rect 23658 33804 23664 33856
rect 23716 33804 23722 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 7006 33600 7012 33652
rect 7064 33640 7070 33652
rect 7064 33612 9352 33640
rect 7064 33600 7070 33612
rect 8570 33532 8576 33584
rect 8628 33532 8634 33584
rect 9324 33572 9352 33612
rect 9490 33600 9496 33652
rect 9548 33600 9554 33652
rect 9858 33600 9864 33652
rect 9916 33640 9922 33652
rect 9953 33643 10011 33649
rect 9953 33640 9965 33643
rect 9916 33612 9965 33640
rect 9916 33600 9922 33612
rect 9953 33609 9965 33612
rect 9999 33609 10011 33643
rect 9953 33603 10011 33609
rect 10226 33600 10232 33652
rect 10284 33640 10290 33652
rect 12253 33643 12311 33649
rect 12253 33640 12265 33643
rect 10284 33612 12265 33640
rect 10284 33600 10290 33612
rect 12253 33609 12265 33612
rect 12299 33609 12311 33643
rect 12253 33603 12311 33609
rect 12713 33643 12771 33649
rect 12713 33609 12725 33643
rect 12759 33640 12771 33643
rect 12802 33640 12808 33652
rect 12759 33612 12808 33640
rect 12759 33609 12771 33612
rect 12713 33603 12771 33609
rect 12802 33600 12808 33612
rect 12860 33600 12866 33652
rect 13906 33600 13912 33652
rect 13964 33600 13970 33652
rect 14918 33600 14924 33652
rect 14976 33640 14982 33652
rect 15105 33643 15163 33649
rect 15105 33640 15117 33643
rect 14976 33612 15117 33640
rect 14976 33600 14982 33612
rect 15105 33609 15117 33612
rect 15151 33609 15163 33643
rect 15105 33603 15163 33609
rect 19521 33643 19579 33649
rect 19521 33609 19533 33643
rect 19567 33640 19579 33643
rect 20714 33640 20720 33652
rect 19567 33612 20720 33640
rect 19567 33609 19579 33612
rect 19521 33603 19579 33609
rect 20714 33600 20720 33612
rect 20772 33600 20778 33652
rect 20806 33600 20812 33652
rect 20864 33640 20870 33652
rect 23842 33640 23848 33652
rect 20864 33612 23848 33640
rect 20864 33600 20870 33612
rect 23842 33600 23848 33612
rect 23900 33600 23906 33652
rect 25225 33643 25283 33649
rect 25225 33640 25237 33643
rect 23952 33612 25237 33640
rect 10321 33575 10379 33581
rect 10321 33572 10333 33575
rect 9324 33544 10333 33572
rect 10321 33541 10333 33544
rect 10367 33541 10379 33575
rect 10321 33535 10379 33541
rect 13817 33575 13875 33581
rect 13817 33541 13829 33575
rect 13863 33572 13875 33575
rect 13998 33572 14004 33584
rect 13863 33544 14004 33572
rect 13863 33541 13875 33544
rect 13817 33535 13875 33541
rect 13998 33532 14004 33544
rect 14056 33572 14062 33584
rect 14734 33572 14740 33584
rect 14056 33544 14740 33572
rect 14056 33532 14062 33544
rect 14734 33532 14740 33544
rect 14792 33532 14798 33584
rect 17126 33572 17132 33584
rect 14936 33544 17132 33572
rect 12621 33507 12679 33513
rect 12621 33473 12633 33507
rect 12667 33504 12679 33507
rect 14936 33504 14964 33544
rect 17126 33532 17132 33544
rect 17184 33532 17190 33584
rect 18601 33575 18659 33581
rect 18601 33541 18613 33575
rect 18647 33572 18659 33575
rect 23290 33572 23296 33584
rect 18647 33544 23296 33572
rect 18647 33541 18659 33544
rect 18601 33535 18659 33541
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 23750 33532 23756 33584
rect 23808 33572 23814 33584
rect 23952 33572 23980 33612
rect 25225 33609 25237 33612
rect 25271 33609 25283 33643
rect 25225 33603 25283 33609
rect 23808 33544 23980 33572
rect 23808 33532 23814 33544
rect 24486 33532 24492 33584
rect 24544 33532 24550 33584
rect 12667 33476 13768 33504
rect 12667 33473 12679 33476
rect 12621 33467 12679 33473
rect 7742 33396 7748 33448
rect 7800 33396 7806 33448
rect 8021 33439 8079 33445
rect 8021 33405 8033 33439
rect 8067 33436 8079 33439
rect 9398 33436 9404 33448
rect 8067 33408 9404 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 9398 33396 9404 33408
rect 9456 33396 9462 33448
rect 10410 33396 10416 33448
rect 10468 33396 10474 33448
rect 10505 33439 10563 33445
rect 10505 33405 10517 33439
rect 10551 33405 10563 33439
rect 10505 33399 10563 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33405 12863 33439
rect 13740 33436 13768 33476
rect 13924 33476 14964 33504
rect 13924 33436 13952 33476
rect 15010 33464 15016 33516
rect 15068 33464 15074 33516
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 18509 33507 18567 33513
rect 15160 33476 18276 33504
rect 15160 33464 15166 33476
rect 13740 33408 13952 33436
rect 14001 33439 14059 33445
rect 12805 33399 12863 33405
rect 14001 33405 14013 33439
rect 14047 33405 14059 33439
rect 14001 33399 14059 33405
rect 10318 33328 10324 33380
rect 10376 33368 10382 33380
rect 10520 33368 10548 33399
rect 10376 33340 10548 33368
rect 10376 33328 10382 33340
rect 11054 33328 11060 33380
rect 11112 33368 11118 33380
rect 12820 33368 12848 33399
rect 11112 33340 12848 33368
rect 11112 33328 11118 33340
rect 13354 33328 13360 33380
rect 13412 33368 13418 33380
rect 14016 33368 14044 33399
rect 14182 33396 14188 33448
rect 14240 33436 14246 33448
rect 15197 33439 15255 33445
rect 15197 33436 15209 33439
rect 14240 33408 15209 33436
rect 14240 33396 14246 33408
rect 15197 33405 15209 33408
rect 15243 33405 15255 33439
rect 15197 33399 15255 33405
rect 18141 33371 18199 33377
rect 18141 33368 18153 33371
rect 13412 33340 14044 33368
rect 14568 33340 18153 33368
rect 13412 33328 13418 33340
rect 10502 33260 10508 33312
rect 10560 33300 10566 33312
rect 12618 33300 12624 33312
rect 10560 33272 12624 33300
rect 10560 33260 10566 33272
rect 12618 33260 12624 33272
rect 12676 33300 12682 33312
rect 13262 33300 13268 33312
rect 12676 33272 13268 33300
rect 12676 33260 12682 33272
rect 13262 33260 13268 33272
rect 13320 33260 13326 33312
rect 13446 33260 13452 33312
rect 13504 33260 13510 33312
rect 13538 33260 13544 33312
rect 13596 33300 13602 33312
rect 14568 33300 14596 33340
rect 18141 33337 18153 33340
rect 18187 33337 18199 33371
rect 18248 33368 18276 33476
rect 18509 33473 18521 33507
rect 18555 33504 18567 33507
rect 18555 33476 18828 33504
rect 18555 33473 18567 33476
rect 18509 33467 18567 33473
rect 18693 33439 18751 33445
rect 18693 33405 18705 33439
rect 18739 33405 18751 33439
rect 18693 33399 18751 33405
rect 18708 33368 18736 33399
rect 18248 33340 18736 33368
rect 18800 33368 18828 33476
rect 18966 33464 18972 33516
rect 19024 33504 19030 33516
rect 19889 33507 19947 33513
rect 19889 33504 19901 33507
rect 19024 33476 19901 33504
rect 19024 33464 19030 33476
rect 19889 33473 19901 33476
rect 19935 33473 19947 33507
rect 21726 33504 21732 33516
rect 19889 33467 19947 33473
rect 20088 33476 21732 33504
rect 19978 33396 19984 33448
rect 20036 33396 20042 33448
rect 20088 33445 20116 33476
rect 21726 33464 21732 33476
rect 21784 33464 21790 33516
rect 20073 33439 20131 33445
rect 20073 33405 20085 33439
rect 20119 33405 20131 33439
rect 20073 33399 20131 33405
rect 20346 33396 20352 33448
rect 20404 33436 20410 33448
rect 22646 33436 22652 33448
rect 20404 33408 22652 33436
rect 20404 33396 20410 33408
rect 22646 33396 22652 33408
rect 22704 33436 22710 33448
rect 23477 33439 23535 33445
rect 23477 33436 23489 33439
rect 22704 33408 23489 33436
rect 22704 33396 22710 33408
rect 23477 33405 23489 33408
rect 23523 33405 23535 33439
rect 23477 33399 23535 33405
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 20162 33368 20168 33380
rect 18800 33340 20168 33368
rect 18141 33331 18199 33337
rect 20162 33328 20168 33340
rect 20220 33328 20226 33380
rect 13596 33272 14596 33300
rect 14645 33303 14703 33309
rect 13596 33260 13602 33272
rect 14645 33269 14657 33303
rect 14691 33300 14703 33303
rect 15102 33300 15108 33312
rect 14691 33272 15108 33300
rect 14691 33269 14703 33272
rect 14645 33263 14703 33269
rect 15102 33260 15108 33272
rect 15160 33260 15166 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 9125 33099 9183 33105
rect 9125 33065 9137 33099
rect 9171 33096 9183 33099
rect 9306 33096 9312 33108
rect 9171 33068 9312 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 9306 33056 9312 33068
rect 9364 33056 9370 33108
rect 9582 33056 9588 33108
rect 9640 33096 9646 33108
rect 11701 33099 11759 33105
rect 11701 33096 11713 33099
rect 9640 33068 11713 33096
rect 9640 33056 9646 33068
rect 11701 33065 11713 33068
rect 11747 33065 11759 33099
rect 11701 33059 11759 33065
rect 12897 33099 12955 33105
rect 12897 33065 12909 33099
rect 12943 33096 12955 33099
rect 15010 33096 15016 33108
rect 12943 33068 15016 33096
rect 12943 33065 12955 33068
rect 12897 33059 12955 33065
rect 15010 33056 15016 33068
rect 15068 33056 15074 33108
rect 18601 33099 18659 33105
rect 18601 33065 18613 33099
rect 18647 33096 18659 33099
rect 20438 33096 20444 33108
rect 18647 33068 20444 33096
rect 18647 33065 18659 33068
rect 18601 33059 18659 33065
rect 20438 33056 20444 33068
rect 20496 33056 20502 33108
rect 20990 33056 20996 33108
rect 21048 33096 21054 33108
rect 21818 33096 21824 33108
rect 21048 33068 21824 33096
rect 21048 33056 21054 33068
rect 21818 33056 21824 33068
rect 21876 33096 21882 33108
rect 22097 33099 22155 33105
rect 22097 33096 22109 33099
rect 21876 33068 22109 33096
rect 21876 33056 21882 33068
rect 22097 33065 22109 33068
rect 22143 33065 22155 33099
rect 22097 33059 22155 33065
rect 23014 33056 23020 33108
rect 23072 33096 23078 33108
rect 23382 33096 23388 33108
rect 23072 33068 23388 33096
rect 23072 33056 23078 33068
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 6822 32988 6828 33040
rect 6880 33028 6886 33040
rect 7285 33031 7343 33037
rect 7285 33028 7297 33031
rect 6880 33000 7297 33028
rect 6880 32988 6886 33000
rect 7285 32997 7297 33000
rect 7331 33028 7343 33031
rect 12710 33028 12716 33040
rect 7331 33000 12716 33028
rect 7331 32997 7343 33000
rect 7285 32991 7343 32997
rect 12710 32988 12716 33000
rect 12768 32988 12774 33040
rect 15838 32988 15844 33040
rect 15896 33028 15902 33040
rect 15896 33000 16988 33028
rect 15896 32988 15902 33000
rect 4890 32920 4896 32972
rect 4948 32960 4954 32972
rect 5537 32963 5595 32969
rect 5537 32960 5549 32963
rect 4948 32932 5549 32960
rect 4948 32920 4954 32932
rect 5537 32929 5549 32932
rect 5583 32960 5595 32963
rect 7742 32960 7748 32972
rect 5583 32932 7748 32960
rect 5583 32929 5595 32932
rect 5537 32923 5595 32929
rect 7742 32920 7748 32932
rect 7800 32920 7806 32972
rect 9398 32920 9404 32972
rect 9456 32960 9462 32972
rect 9677 32963 9735 32969
rect 9677 32960 9689 32963
rect 9456 32932 9689 32960
rect 9456 32920 9462 32932
rect 9677 32929 9689 32932
rect 9723 32929 9735 32963
rect 12253 32963 12311 32969
rect 12253 32960 12265 32963
rect 9677 32923 9735 32929
rect 9784 32932 12265 32960
rect 8386 32852 8392 32904
rect 8444 32892 8450 32904
rect 9784 32892 9812 32932
rect 12253 32929 12265 32932
rect 12299 32929 12311 32963
rect 12253 32923 12311 32929
rect 13541 32963 13599 32969
rect 13541 32929 13553 32963
rect 13587 32960 13599 32963
rect 13814 32960 13820 32972
rect 13587 32932 13820 32960
rect 13587 32929 13599 32932
rect 13541 32923 13599 32929
rect 13814 32920 13820 32932
rect 13872 32920 13878 32972
rect 16114 32920 16120 32972
rect 16172 32920 16178 32972
rect 16298 32920 16304 32972
rect 16356 32920 16362 32972
rect 16850 32920 16856 32972
rect 16908 32920 16914 32972
rect 16960 32960 16988 33000
rect 18966 32988 18972 33040
rect 19024 33028 19030 33040
rect 19610 33028 19616 33040
rect 19024 33000 19616 33028
rect 19024 32988 19030 33000
rect 19610 32988 19616 33000
rect 19668 32988 19674 33040
rect 16960 32932 18368 32960
rect 8444 32864 9812 32892
rect 12069 32895 12127 32901
rect 8444 32852 8450 32864
rect 12069 32861 12081 32895
rect 12115 32892 12127 32895
rect 12158 32892 12164 32904
rect 12115 32864 12164 32892
rect 12115 32861 12127 32864
rect 12069 32855 12127 32861
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 13357 32895 13415 32901
rect 13357 32861 13369 32895
rect 13403 32892 13415 32895
rect 13630 32892 13636 32904
rect 13403 32864 13636 32892
rect 13403 32861 13415 32864
rect 13357 32855 13415 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 16025 32895 16083 32901
rect 16025 32861 16037 32895
rect 16071 32892 16083 32895
rect 16574 32892 16580 32904
rect 16071 32864 16580 32892
rect 16071 32861 16083 32864
rect 16025 32855 16083 32861
rect 16574 32852 16580 32864
rect 16632 32852 16638 32904
rect 5813 32827 5871 32833
rect 5813 32793 5825 32827
rect 5859 32793 5871 32827
rect 5813 32787 5871 32793
rect 5828 32756 5856 32787
rect 6546 32784 6552 32836
rect 6604 32784 6610 32836
rect 8662 32784 8668 32836
rect 8720 32824 8726 32836
rect 9493 32827 9551 32833
rect 9493 32824 9505 32827
rect 8720 32796 9505 32824
rect 8720 32784 8726 32796
rect 9493 32793 9505 32796
rect 9539 32793 9551 32827
rect 9493 32787 9551 32793
rect 16206 32784 16212 32836
rect 16264 32824 16270 32836
rect 17129 32827 17187 32833
rect 17129 32824 17141 32827
rect 16264 32796 17141 32824
rect 16264 32784 16270 32796
rect 17129 32793 17141 32796
rect 17175 32793 17187 32827
rect 18340 32824 18368 32932
rect 20346 32920 20352 32972
rect 20404 32920 20410 32972
rect 20625 32963 20683 32969
rect 20625 32929 20637 32963
rect 20671 32960 20683 32963
rect 22462 32960 22468 32972
rect 20671 32932 22468 32960
rect 20671 32929 20683 32932
rect 20625 32923 20683 32929
rect 22462 32920 22468 32932
rect 22520 32960 22526 32972
rect 23106 32960 23112 32972
rect 22520 32932 23112 32960
rect 22520 32920 22526 32932
rect 23106 32920 23112 32932
rect 23164 32920 23170 32972
rect 23201 32963 23259 32969
rect 23201 32929 23213 32963
rect 23247 32960 23259 32963
rect 23382 32960 23388 32972
rect 23247 32932 23388 32960
rect 23247 32929 23259 32932
rect 23201 32923 23259 32929
rect 23382 32920 23388 32932
rect 23440 32920 23446 32972
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19705 32895 19763 32901
rect 19705 32892 19717 32895
rect 19208 32864 19717 32892
rect 19208 32852 19214 32864
rect 19705 32861 19717 32864
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 22925 32895 22983 32901
rect 22925 32861 22937 32895
rect 22971 32892 22983 32895
rect 23290 32892 23296 32904
rect 22971 32864 23296 32892
rect 22971 32861 22983 32864
rect 22925 32855 22983 32861
rect 23290 32852 23296 32864
rect 23348 32852 23354 32904
rect 24029 32895 24087 32901
rect 24029 32861 24041 32895
rect 24075 32892 24087 32895
rect 24854 32892 24860 32904
rect 24075 32864 24860 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 25314 32852 25320 32904
rect 25372 32852 25378 32904
rect 19058 32824 19064 32836
rect 18340 32810 19064 32824
rect 18354 32796 19064 32810
rect 17129 32787 17187 32793
rect 19058 32784 19064 32796
rect 19116 32784 19122 32836
rect 20714 32824 20720 32836
rect 19444 32796 20720 32824
rect 6822 32756 6828 32768
rect 5828 32728 6828 32756
rect 6822 32716 6828 32728
rect 6880 32716 6886 32768
rect 9306 32716 9312 32768
rect 9364 32756 9370 32768
rect 9585 32759 9643 32765
rect 9585 32756 9597 32759
rect 9364 32728 9597 32756
rect 9364 32716 9370 32728
rect 9585 32725 9597 32728
rect 9631 32725 9643 32759
rect 9585 32719 9643 32725
rect 12066 32716 12072 32768
rect 12124 32756 12130 32768
rect 12161 32759 12219 32765
rect 12161 32756 12173 32759
rect 12124 32728 12173 32756
rect 12124 32716 12130 32728
rect 12161 32725 12173 32728
rect 12207 32725 12219 32759
rect 12161 32719 12219 32725
rect 13262 32716 13268 32768
rect 13320 32716 13326 32768
rect 14734 32716 14740 32768
rect 14792 32756 14798 32768
rect 15657 32759 15715 32765
rect 15657 32756 15669 32759
rect 14792 32728 15669 32756
rect 14792 32716 14798 32728
rect 15657 32725 15669 32728
rect 15703 32725 15715 32759
rect 15657 32719 15715 32725
rect 17034 32716 17040 32768
rect 17092 32756 17098 32768
rect 19444 32756 19472 32796
rect 20714 32784 20720 32796
rect 20772 32784 20778 32836
rect 21910 32824 21916 32836
rect 21850 32796 21916 32824
rect 21910 32784 21916 32796
rect 21968 32784 21974 32836
rect 23014 32784 23020 32836
rect 23072 32784 23078 32836
rect 17092 32728 19472 32756
rect 19521 32759 19579 32765
rect 17092 32716 17098 32728
rect 19521 32725 19533 32759
rect 19567 32756 19579 32759
rect 21542 32756 21548 32768
rect 19567 32728 21548 32756
rect 19567 32725 19579 32728
rect 19521 32719 19579 32725
rect 21542 32716 21548 32728
rect 21600 32716 21606 32768
rect 22554 32716 22560 32768
rect 22612 32716 22618 32768
rect 23566 32716 23572 32768
rect 23624 32756 23630 32768
rect 23845 32759 23903 32765
rect 23845 32756 23857 32759
rect 23624 32728 23857 32756
rect 23624 32716 23630 32728
rect 23845 32725 23857 32728
rect 23891 32725 23903 32759
rect 23845 32719 23903 32725
rect 25130 32716 25136 32768
rect 25188 32716 25194 32768
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 8570 32512 8576 32564
rect 8628 32552 8634 32564
rect 14826 32552 14832 32564
rect 8628 32524 10548 32552
rect 8628 32512 8634 32524
rect 9401 32487 9459 32493
rect 9401 32453 9413 32487
rect 9447 32484 9459 32487
rect 9490 32484 9496 32496
rect 9447 32456 9496 32484
rect 9447 32453 9459 32456
rect 9401 32447 9459 32453
rect 9490 32444 9496 32456
rect 9548 32444 9554 32496
rect 10520 32428 10548 32524
rect 10888 32524 14832 32552
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1765 32419 1823 32425
rect 1765 32416 1777 32419
rect 992 32388 1777 32416
rect 992 32376 998 32388
rect 1765 32385 1777 32388
rect 1811 32385 1823 32419
rect 1765 32379 1823 32385
rect 7742 32376 7748 32428
rect 7800 32416 7806 32428
rect 9125 32419 9183 32425
rect 9125 32416 9137 32419
rect 7800 32388 9137 32416
rect 7800 32376 7806 32388
rect 9125 32385 9137 32388
rect 9171 32385 9183 32419
rect 9125 32379 9183 32385
rect 10502 32376 10508 32428
rect 10560 32376 10566 32428
rect 8662 32308 8668 32360
rect 8720 32308 8726 32360
rect 1578 32172 1584 32224
rect 1636 32172 1642 32224
rect 7650 32172 7656 32224
rect 7708 32172 7714 32224
rect 9766 32172 9772 32224
rect 9824 32212 9830 32224
rect 10888 32221 10916 32524
rect 14826 32512 14832 32524
rect 14884 32512 14890 32564
rect 17310 32512 17316 32564
rect 17368 32512 17374 32564
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 19429 32555 19487 32561
rect 19429 32552 19441 32555
rect 19392 32524 19441 32552
rect 19392 32512 19398 32524
rect 19429 32521 19441 32524
rect 19475 32521 19487 32555
rect 19429 32515 19487 32521
rect 19521 32555 19579 32561
rect 19521 32521 19533 32555
rect 19567 32552 19579 32555
rect 19702 32552 19708 32564
rect 19567 32524 19708 32552
rect 19567 32521 19579 32524
rect 19521 32515 19579 32521
rect 19702 32512 19708 32524
rect 19760 32512 19766 32564
rect 20901 32555 20959 32561
rect 20901 32521 20913 32555
rect 20947 32552 20959 32555
rect 21266 32552 21272 32564
rect 20947 32524 21272 32552
rect 20947 32521 20959 32524
rect 20901 32515 20959 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 22278 32512 22284 32564
rect 22336 32552 22342 32564
rect 23109 32555 23167 32561
rect 23109 32552 23121 32555
rect 22336 32524 23121 32552
rect 22336 32512 22342 32524
rect 23109 32521 23121 32524
rect 23155 32552 23167 32555
rect 25130 32552 25136 32564
rect 23155 32524 25136 32552
rect 23155 32521 23167 32524
rect 23109 32515 23167 32521
rect 25130 32512 25136 32524
rect 25188 32512 25194 32564
rect 16758 32444 16764 32496
rect 16816 32484 16822 32496
rect 17221 32487 17279 32493
rect 17221 32484 17233 32487
rect 16816 32456 17233 32484
rect 16816 32444 16822 32456
rect 17221 32453 17233 32456
rect 17267 32453 17279 32487
rect 17221 32447 17279 32453
rect 17402 32444 17408 32496
rect 17460 32484 17466 32496
rect 20806 32484 20812 32496
rect 17460 32456 20812 32484
rect 17460 32444 17466 32456
rect 20806 32444 20812 32456
rect 20864 32444 20870 32496
rect 20993 32487 21051 32493
rect 20993 32453 21005 32487
rect 21039 32484 21051 32487
rect 21358 32484 21364 32496
rect 21039 32456 21364 32484
rect 21039 32453 21051 32456
rect 20993 32447 21051 32453
rect 21358 32444 21364 32456
rect 21416 32444 21422 32496
rect 21836 32456 24072 32484
rect 13262 32376 13268 32428
rect 13320 32416 13326 32428
rect 13449 32419 13507 32425
rect 13449 32416 13461 32419
rect 13320 32388 13461 32416
rect 13320 32376 13326 32388
rect 13449 32385 13461 32388
rect 13495 32385 13507 32419
rect 13449 32379 13507 32385
rect 15838 32376 15844 32428
rect 15896 32376 15902 32428
rect 18414 32416 18420 32428
rect 17420 32388 18420 32416
rect 14458 32308 14464 32360
rect 14516 32308 14522 32360
rect 14737 32351 14795 32357
rect 14737 32317 14749 32351
rect 14783 32348 14795 32351
rect 16758 32348 16764 32360
rect 14783 32320 16764 32348
rect 14783 32317 14795 32320
rect 14737 32311 14795 32317
rect 16758 32308 16764 32320
rect 16816 32348 16822 32360
rect 17420 32348 17448 32388
rect 18414 32376 18420 32388
rect 18472 32376 18478 32428
rect 20254 32376 20260 32428
rect 20312 32416 20318 32428
rect 21836 32416 21864 32456
rect 20312 32388 21864 32416
rect 20312 32376 20318 32388
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 23017 32419 23075 32425
rect 23017 32385 23029 32419
rect 23063 32416 23075 32419
rect 23290 32416 23296 32428
rect 23063 32388 23296 32416
rect 23063 32385 23075 32388
rect 23017 32379 23075 32385
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 24044 32425 24072 32456
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 16816 32320 17448 32348
rect 17497 32351 17555 32357
rect 16816 32308 16822 32320
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 18966 32348 18972 32360
rect 17543 32320 18972 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 18966 32308 18972 32320
rect 19024 32308 19030 32360
rect 19613 32351 19671 32357
rect 19613 32317 19625 32351
rect 19659 32317 19671 32351
rect 19613 32311 19671 32317
rect 17034 32240 17040 32292
rect 17092 32280 17098 32292
rect 17402 32280 17408 32292
rect 17092 32252 17408 32280
rect 17092 32240 17098 32252
rect 17402 32240 17408 32252
rect 17460 32240 17466 32292
rect 17586 32240 17592 32292
rect 17644 32280 17650 32292
rect 19628 32280 19656 32311
rect 20806 32308 20812 32360
rect 20864 32348 20870 32360
rect 21085 32351 21143 32357
rect 21085 32348 21097 32351
rect 20864 32320 21097 32348
rect 20864 32308 20870 32320
rect 21085 32317 21097 32320
rect 21131 32317 21143 32351
rect 21085 32311 21143 32317
rect 23198 32308 23204 32360
rect 23256 32308 23262 32360
rect 17644 32252 19656 32280
rect 17644 32240 17650 32252
rect 20990 32240 20996 32292
rect 21048 32280 21054 32292
rect 25133 32283 25191 32289
rect 25133 32280 25145 32283
rect 21048 32252 25145 32280
rect 21048 32240 21054 32252
rect 25133 32249 25145 32252
rect 25179 32249 25191 32283
rect 25133 32243 25191 32249
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 9824 32184 10885 32212
rect 9824 32172 9830 32184
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 10873 32175 10931 32181
rect 12342 32172 12348 32224
rect 12400 32212 12406 32224
rect 14274 32212 14280 32224
rect 12400 32184 14280 32212
rect 12400 32172 12406 32184
rect 14274 32172 14280 32184
rect 14332 32172 14338 32224
rect 14550 32172 14556 32224
rect 14608 32212 14614 32224
rect 16209 32215 16267 32221
rect 16209 32212 16221 32215
rect 14608 32184 16221 32212
rect 14608 32172 14614 32184
rect 16209 32181 16221 32184
rect 16255 32212 16267 32215
rect 16298 32212 16304 32224
rect 16255 32184 16304 32212
rect 16255 32181 16267 32184
rect 16209 32175 16267 32181
rect 16298 32172 16304 32184
rect 16356 32172 16362 32224
rect 16853 32215 16911 32221
rect 16853 32181 16865 32215
rect 16899 32212 16911 32215
rect 17770 32212 17776 32224
rect 16899 32184 17776 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 17770 32172 17776 32184
rect 17828 32172 17834 32224
rect 18414 32172 18420 32224
rect 18472 32212 18478 32224
rect 19061 32215 19119 32221
rect 19061 32212 19073 32215
rect 18472 32184 19073 32212
rect 18472 32172 18478 32184
rect 19061 32181 19073 32184
rect 19107 32181 19119 32215
rect 19061 32175 19119 32181
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 20438 32212 20444 32224
rect 19392 32184 20444 32212
rect 19392 32172 19398 32184
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 20530 32172 20536 32224
rect 20588 32172 20594 32224
rect 22002 32172 22008 32224
rect 22060 32172 22066 32224
rect 22186 32172 22192 32224
rect 22244 32212 22250 32224
rect 22649 32215 22707 32221
rect 22649 32212 22661 32215
rect 22244 32184 22661 32212
rect 22244 32172 22250 32184
rect 22649 32181 22661 32184
rect 22695 32181 22707 32215
rect 22649 32175 22707 32181
rect 22830 32172 22836 32224
rect 22888 32212 22894 32224
rect 23474 32212 23480 32224
rect 22888 32184 23480 32212
rect 22888 32172 22894 32184
rect 23474 32172 23480 32184
rect 23532 32172 23538 32224
rect 23845 32215 23903 32221
rect 23845 32181 23857 32215
rect 23891 32212 23903 32215
rect 24302 32212 24308 32224
rect 23891 32184 24308 32212
rect 23891 32181 23903 32184
rect 23845 32175 23903 32181
rect 24302 32172 24308 32184
rect 24360 32172 24366 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 6914 31968 6920 32020
rect 6972 31968 6978 32020
rect 7469 32011 7527 32017
rect 7469 31977 7481 32011
rect 7515 32008 7527 32011
rect 7834 32008 7840 32020
rect 7515 31980 7840 32008
rect 7515 31977 7527 31980
rect 7469 31971 7527 31977
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 9398 31968 9404 32020
rect 9456 32008 9462 32020
rect 10873 32011 10931 32017
rect 10873 32008 10885 32011
rect 9456 31980 10885 32008
rect 9456 31968 9462 31980
rect 10873 31977 10885 31980
rect 10919 32008 10931 32011
rect 11054 32008 11060 32020
rect 10919 31980 11060 32008
rect 10919 31977 10931 31980
rect 10873 31971 10931 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 11974 31968 11980 32020
rect 12032 32008 12038 32020
rect 12345 32011 12403 32017
rect 12345 32008 12357 32011
rect 12032 31980 12357 32008
rect 12032 31968 12038 31980
rect 12345 31977 12357 31980
rect 12391 31977 12403 32011
rect 19978 32008 19984 32020
rect 12345 31971 12403 31977
rect 14384 31980 19984 32008
rect 4890 31832 4896 31884
rect 4948 31872 4954 31884
rect 5169 31875 5227 31881
rect 5169 31872 5181 31875
rect 4948 31844 5181 31872
rect 4948 31832 4954 31844
rect 5169 31841 5181 31844
rect 5215 31841 5227 31875
rect 5169 31835 5227 31841
rect 5445 31875 5503 31881
rect 5445 31841 5457 31875
rect 5491 31872 5503 31875
rect 8113 31875 8171 31881
rect 8113 31872 8125 31875
rect 5491 31844 8125 31872
rect 5491 31841 5503 31844
rect 5445 31835 5503 31841
rect 8113 31841 8125 31844
rect 8159 31872 8171 31875
rect 8386 31872 8392 31884
rect 8159 31844 8392 31872
rect 8159 31841 8171 31844
rect 8113 31835 8171 31841
rect 8386 31832 8392 31844
rect 8444 31832 8450 31884
rect 8478 31832 8484 31884
rect 8536 31872 8542 31884
rect 9401 31875 9459 31881
rect 9401 31872 9413 31875
rect 8536 31844 9413 31872
rect 8536 31832 8542 31844
rect 9401 31841 9413 31844
rect 9447 31872 9459 31875
rect 9490 31872 9496 31884
rect 9447 31844 9496 31872
rect 9447 31841 9459 31844
rect 9401 31835 9459 31841
rect 9490 31832 9496 31844
rect 9548 31872 9554 31884
rect 9548 31844 11008 31872
rect 9548 31832 9554 31844
rect 4706 31764 4712 31816
rect 4764 31764 4770 31816
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 7929 31807 7987 31813
rect 7929 31773 7941 31807
rect 7975 31804 7987 31807
rect 8938 31804 8944 31816
rect 7975 31776 8944 31804
rect 7975 31773 7987 31776
rect 7929 31767 7987 31773
rect 8938 31764 8944 31776
rect 8996 31764 9002 31816
rect 9122 31764 9128 31816
rect 9180 31764 9186 31816
rect 10502 31764 10508 31816
rect 10560 31764 10566 31816
rect 7834 31628 7840 31680
rect 7892 31628 7898 31680
rect 10318 31628 10324 31680
rect 10376 31668 10382 31680
rect 10520 31668 10548 31764
rect 10980 31736 11008 31844
rect 12710 31832 12716 31884
rect 12768 31872 12774 31884
rect 12897 31875 12955 31881
rect 12897 31872 12909 31875
rect 12768 31844 12909 31872
rect 12768 31832 12774 31844
rect 12897 31841 12909 31844
rect 12943 31841 12955 31875
rect 12897 31835 12955 31841
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31804 12863 31807
rect 14384 31804 14412 31980
rect 19978 31968 19984 31980
rect 20036 32008 20042 32020
rect 20346 32008 20352 32020
rect 20036 31980 20352 32008
rect 20036 31968 20042 31980
rect 20346 31968 20352 31980
rect 20404 31968 20410 32020
rect 21358 31968 21364 32020
rect 21416 32008 21422 32020
rect 23845 32011 23903 32017
rect 23845 32008 23857 32011
rect 21416 31980 23857 32008
rect 21416 31968 21422 31980
rect 23845 31977 23857 31980
rect 23891 31977 23903 32011
rect 23845 31971 23903 31977
rect 16482 31900 16488 31952
rect 16540 31940 16546 31952
rect 16540 31912 17172 31940
rect 16540 31900 16546 31912
rect 14458 31832 14464 31884
rect 14516 31872 14522 31884
rect 15105 31875 15163 31881
rect 15105 31872 15117 31875
rect 14516 31844 15117 31872
rect 14516 31832 14522 31844
rect 15105 31841 15117 31844
rect 15151 31872 15163 31875
rect 16850 31872 16856 31884
rect 15151 31844 16856 31872
rect 15151 31841 15163 31844
rect 15105 31835 15163 31841
rect 16850 31832 16856 31844
rect 16908 31832 16914 31884
rect 12851 31776 14412 31804
rect 17144 31804 17172 31912
rect 17218 31900 17224 31952
rect 17276 31940 17282 31952
rect 17313 31943 17371 31949
rect 17313 31940 17325 31943
rect 17276 31912 17325 31940
rect 17276 31900 17282 31912
rect 17313 31909 17325 31912
rect 17359 31909 17371 31943
rect 17313 31903 17371 31909
rect 17494 31900 17500 31952
rect 17552 31940 17558 31952
rect 19429 31943 19487 31949
rect 17552 31912 18000 31940
rect 17552 31900 17558 31912
rect 17770 31832 17776 31884
rect 17828 31832 17834 31884
rect 17862 31832 17868 31884
rect 17920 31832 17926 31884
rect 17972 31872 18000 31912
rect 19429 31909 19441 31943
rect 19475 31940 19487 31943
rect 20438 31940 20444 31952
rect 19475 31912 20444 31940
rect 19475 31909 19487 31912
rect 19429 31903 19487 31909
rect 20438 31900 20444 31912
rect 20496 31900 20502 31952
rect 20625 31943 20683 31949
rect 20625 31909 20637 31943
rect 20671 31940 20683 31943
rect 21726 31940 21732 31952
rect 20671 31912 21732 31940
rect 20671 31909 20683 31912
rect 20625 31903 20683 31909
rect 21726 31900 21732 31912
rect 21784 31900 21790 31952
rect 21821 31943 21879 31949
rect 21821 31909 21833 31943
rect 21867 31940 21879 31943
rect 22278 31940 22284 31952
rect 21867 31912 22284 31940
rect 21867 31909 21879 31912
rect 21821 31903 21879 31909
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 23201 31943 23259 31949
rect 23201 31909 23213 31943
rect 23247 31940 23259 31943
rect 23290 31940 23296 31952
rect 23247 31912 23296 31940
rect 23247 31909 23259 31912
rect 23201 31903 23259 31909
rect 23290 31900 23296 31912
rect 23348 31900 23354 31952
rect 24581 31943 24639 31949
rect 24581 31909 24593 31943
rect 24627 31940 24639 31943
rect 24670 31940 24676 31952
rect 24627 31912 24676 31940
rect 24627 31909 24639 31912
rect 24581 31903 24639 31909
rect 24670 31900 24676 31912
rect 24728 31900 24734 31952
rect 20990 31872 20996 31884
rect 17972 31844 20996 31872
rect 20990 31832 20996 31844
rect 21048 31832 21054 31884
rect 21082 31832 21088 31884
rect 21140 31872 21146 31884
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 21140 31844 21189 31872
rect 21140 31832 21146 31844
rect 21177 31841 21189 31844
rect 21223 31872 21235 31875
rect 22465 31875 22523 31881
rect 22465 31872 22477 31875
rect 21223 31844 22477 31872
rect 21223 31841 21235 31844
rect 21177 31835 21235 31841
rect 22465 31841 22477 31844
rect 22511 31872 22523 31875
rect 23014 31872 23020 31884
rect 22511 31844 23020 31872
rect 22511 31841 22523 31844
rect 22465 31835 22523 31841
rect 23014 31832 23020 31844
rect 23072 31832 23078 31884
rect 23474 31832 23480 31884
rect 23532 31872 23538 31884
rect 23532 31844 24808 31872
rect 23532 31832 23538 31844
rect 19613 31807 19671 31813
rect 19613 31804 19625 31807
rect 17144 31776 19625 31804
rect 12851 31773 12863 31776
rect 12805 31767 12863 31773
rect 19613 31773 19625 31776
rect 19659 31773 19671 31807
rect 21910 31804 21916 31816
rect 19613 31767 19671 31773
rect 21008 31776 21916 31804
rect 15286 31736 15292 31748
rect 10980 31708 15292 31736
rect 15286 31696 15292 31708
rect 15344 31696 15350 31748
rect 15378 31696 15384 31748
rect 15436 31696 15442 31748
rect 15838 31736 15844 31748
rect 15488 31708 15844 31736
rect 10376 31640 10548 31668
rect 10376 31628 10382 31640
rect 12710 31628 12716 31680
rect 12768 31628 12774 31680
rect 15194 31628 15200 31680
rect 15252 31668 15258 31680
rect 15488 31668 15516 31708
rect 15838 31696 15844 31708
rect 15896 31696 15902 31748
rect 17681 31739 17739 31745
rect 17681 31705 17693 31739
rect 17727 31736 17739 31739
rect 18690 31736 18696 31748
rect 17727 31708 18696 31736
rect 17727 31705 17739 31708
rect 17681 31699 17739 31705
rect 18690 31696 18696 31708
rect 18748 31696 18754 31748
rect 20622 31696 20628 31748
rect 20680 31736 20686 31748
rect 21008 31745 21036 31776
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 24026 31764 24032 31816
rect 24084 31764 24090 31816
rect 24780 31813 24808 31844
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 20993 31739 21051 31745
rect 20993 31736 21005 31739
rect 20680 31708 21005 31736
rect 20680 31696 20686 31708
rect 20993 31705 21005 31708
rect 21039 31705 21051 31739
rect 20993 31699 21051 31705
rect 21085 31739 21143 31745
rect 21085 31705 21097 31739
rect 21131 31736 21143 31739
rect 21450 31736 21456 31748
rect 21131 31708 21456 31736
rect 21131 31705 21143 31708
rect 21085 31699 21143 31705
rect 21450 31696 21456 31708
rect 21508 31696 21514 31748
rect 22189 31739 22247 31745
rect 22189 31705 22201 31739
rect 22235 31736 22247 31739
rect 25590 31736 25596 31748
rect 22235 31708 25596 31736
rect 22235 31705 22247 31708
rect 22189 31699 22247 31705
rect 15252 31640 15516 31668
rect 15252 31628 15258 31640
rect 16758 31628 16764 31680
rect 16816 31668 16822 31680
rect 16853 31671 16911 31677
rect 16853 31668 16865 31671
rect 16816 31640 16865 31668
rect 16816 31628 16822 31640
rect 16853 31637 16865 31640
rect 16899 31637 16911 31671
rect 16853 31631 16911 31637
rect 19702 31628 19708 31680
rect 19760 31668 19766 31680
rect 20070 31668 20076 31680
rect 19760 31640 20076 31668
rect 19760 31628 19766 31640
rect 20070 31628 20076 31640
rect 20128 31668 20134 31680
rect 22204 31668 22232 31699
rect 25590 31696 25596 31708
rect 25648 31696 25654 31748
rect 20128 31640 22232 31668
rect 22281 31671 22339 31677
rect 20128 31628 20134 31640
rect 22281 31637 22293 31671
rect 22327 31668 22339 31671
rect 22922 31668 22928 31680
rect 22327 31640 22928 31668
rect 22327 31637 22339 31640
rect 22281 31631 22339 31637
rect 22922 31628 22928 31640
rect 22980 31628 22986 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 4525 31467 4583 31473
rect 4525 31433 4537 31467
rect 4571 31464 4583 31467
rect 4614 31464 4620 31476
rect 4571 31436 4620 31464
rect 4571 31433 4583 31436
rect 4525 31427 4583 31433
rect 4614 31424 4620 31436
rect 4672 31424 4678 31476
rect 4706 31424 4712 31476
rect 4764 31464 4770 31476
rect 4893 31467 4951 31473
rect 4893 31464 4905 31467
rect 4764 31436 4905 31464
rect 4764 31424 4770 31436
rect 4893 31433 4905 31436
rect 4939 31433 4951 31467
rect 4893 31427 4951 31433
rect 7006 31424 7012 31476
rect 7064 31424 7070 31476
rect 10042 31424 10048 31476
rect 10100 31464 10106 31476
rect 10137 31467 10195 31473
rect 10137 31464 10149 31467
rect 10100 31436 10149 31464
rect 10100 31424 10106 31436
rect 10137 31433 10149 31436
rect 10183 31433 10195 31467
rect 10137 31427 10195 31433
rect 10597 31467 10655 31473
rect 10597 31433 10609 31467
rect 10643 31464 10655 31467
rect 10778 31464 10784 31476
rect 10643 31436 10784 31464
rect 10643 31433 10655 31436
rect 10597 31427 10655 31433
rect 10778 31424 10784 31436
rect 10836 31424 10842 31476
rect 17126 31424 17132 31476
rect 17184 31464 17190 31476
rect 17313 31467 17371 31473
rect 17313 31464 17325 31467
rect 17184 31436 17325 31464
rect 17184 31424 17190 31436
rect 17313 31433 17325 31436
rect 17359 31433 17371 31467
rect 17313 31427 17371 31433
rect 4985 31399 5043 31405
rect 4985 31365 4997 31399
rect 5031 31396 5043 31399
rect 5074 31396 5080 31408
rect 5031 31368 5080 31396
rect 5031 31365 5043 31368
rect 4985 31359 5043 31365
rect 5074 31356 5080 31368
rect 5132 31356 5138 31408
rect 19426 31356 19432 31408
rect 19484 31396 19490 31408
rect 24857 31399 24915 31405
rect 19484 31368 22094 31396
rect 19484 31356 19490 31368
rect 4154 31288 4160 31340
rect 4212 31328 4218 31340
rect 4212 31300 6914 31328
rect 4212 31288 4218 31300
rect 5169 31263 5227 31269
rect 5169 31229 5181 31263
rect 5215 31260 5227 31263
rect 5350 31260 5356 31272
rect 5215 31232 5356 31260
rect 5215 31229 5227 31232
rect 5169 31223 5227 31229
rect 5350 31220 5356 31232
rect 5408 31220 5414 31272
rect 6886 31260 6914 31300
rect 7374 31288 7380 31340
rect 7432 31288 7438 31340
rect 7834 31288 7840 31340
rect 7892 31328 7898 31340
rect 8389 31331 8447 31337
rect 8389 31328 8401 31331
rect 7892 31300 8401 31328
rect 7892 31288 7898 31300
rect 8389 31297 8401 31300
rect 8435 31297 8447 31331
rect 8389 31291 8447 31297
rect 10505 31331 10563 31337
rect 10505 31297 10517 31331
rect 10551 31297 10563 31331
rect 10505 31291 10563 31297
rect 7466 31260 7472 31272
rect 6886 31232 7472 31260
rect 7466 31220 7472 31232
rect 7524 31220 7530 31272
rect 7558 31220 7564 31272
rect 7616 31220 7622 31272
rect 10520 31204 10548 31291
rect 17678 31288 17684 31340
rect 17736 31288 17742 31340
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31328 17831 31331
rect 20806 31328 20812 31340
rect 17819 31300 20812 31328
rect 17819 31297 17831 31300
rect 17773 31291 17831 31297
rect 20806 31288 20812 31300
rect 20864 31288 20870 31340
rect 22066 31328 22094 31368
rect 24857 31365 24869 31399
rect 24903 31396 24915 31399
rect 25866 31396 25872 31408
rect 24903 31368 25872 31396
rect 24903 31365 24915 31368
rect 24857 31359 24915 31365
rect 25866 31356 25872 31368
rect 25924 31356 25930 31408
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 22066 31300 22201 31328
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22189 31291 22247 31297
rect 22830 31288 22836 31340
rect 22888 31328 22894 31340
rect 23569 31331 23627 31337
rect 23569 31328 23581 31331
rect 22888 31300 23581 31328
rect 22888 31288 22894 31300
rect 23569 31297 23581 31300
rect 23615 31297 23627 31331
rect 23569 31291 23627 31297
rect 24394 31288 24400 31340
rect 24452 31328 24458 31340
rect 24673 31331 24731 31337
rect 24673 31328 24685 31331
rect 24452 31300 24685 31328
rect 24452 31288 24458 31300
rect 24673 31297 24685 31300
rect 24719 31297 24731 31331
rect 24673 31291 24731 31297
rect 10686 31220 10692 31272
rect 10744 31220 10750 31272
rect 15286 31220 15292 31272
rect 15344 31260 15350 31272
rect 17865 31263 17923 31269
rect 17865 31260 17877 31263
rect 15344 31232 17877 31260
rect 15344 31220 15350 31232
rect 17865 31229 17877 31232
rect 17911 31229 17923 31263
rect 17865 31223 17923 31229
rect 5442 31152 5448 31204
rect 5500 31192 5506 31204
rect 10502 31192 10508 31204
rect 5500 31164 10508 31192
rect 5500 31152 5506 31164
rect 10502 31152 10508 31164
rect 10560 31152 10566 31204
rect 18782 31152 18788 31204
rect 18840 31192 18846 31204
rect 21450 31192 21456 31204
rect 18840 31164 21456 31192
rect 18840 31152 18846 31164
rect 21450 31152 21456 31164
rect 21508 31152 21514 31204
rect 22005 31195 22063 31201
rect 22005 31161 22017 31195
rect 22051 31192 22063 31195
rect 25222 31192 25228 31204
rect 22051 31164 25228 31192
rect 22051 31161 22063 31164
rect 22005 31155 22063 31161
rect 25222 31152 25228 31164
rect 25280 31152 25286 31204
rect 23385 31127 23443 31133
rect 23385 31093 23397 31127
rect 23431 31124 23443 31127
rect 23842 31124 23848 31136
rect 23431 31096 23848 31124
rect 23431 31093 23443 31096
rect 23385 31087 23443 31093
rect 23842 31084 23848 31096
rect 23900 31084 23906 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 7374 30880 7380 30932
rect 7432 30920 7438 30932
rect 8389 30923 8447 30929
rect 8389 30920 8401 30923
rect 7432 30892 8401 30920
rect 7432 30880 7438 30892
rect 8389 30889 8401 30892
rect 8435 30889 8447 30923
rect 8389 30883 8447 30889
rect 11044 30923 11102 30929
rect 11044 30889 11056 30923
rect 11090 30920 11102 30923
rect 11238 30920 11244 30932
rect 11090 30892 11244 30920
rect 11090 30889 11102 30892
rect 11044 30883 11102 30889
rect 11238 30880 11244 30892
rect 11296 30920 11302 30932
rect 13354 30920 13360 30932
rect 11296 30892 13360 30920
rect 11296 30880 11302 30892
rect 13354 30880 13360 30892
rect 13412 30880 13418 30932
rect 7009 30855 7067 30861
rect 7009 30821 7021 30855
rect 7055 30852 7067 30855
rect 7742 30852 7748 30864
rect 7055 30824 7748 30852
rect 7055 30821 7067 30824
rect 7009 30815 7067 30821
rect 7742 30812 7748 30824
rect 7800 30812 7806 30864
rect 12250 30812 12256 30864
rect 12308 30852 12314 30864
rect 12989 30855 13047 30861
rect 12989 30852 13001 30855
rect 12308 30824 13001 30852
rect 12308 30812 12314 30824
rect 12989 30821 13001 30824
rect 13035 30821 13047 30855
rect 12989 30815 13047 30821
rect 13464 30824 14320 30852
rect 6270 30744 6276 30796
rect 6328 30784 6334 30796
rect 7190 30784 7196 30796
rect 6328 30756 7196 30784
rect 6328 30744 6334 30756
rect 7190 30744 7196 30756
rect 7248 30784 7254 30796
rect 7469 30787 7527 30793
rect 7469 30784 7481 30787
rect 7248 30756 7481 30784
rect 7248 30744 7254 30756
rect 7469 30753 7481 30756
rect 7515 30753 7527 30787
rect 7469 30747 7527 30753
rect 7561 30787 7619 30793
rect 7561 30753 7573 30787
rect 7607 30784 7619 30787
rect 7607 30756 9076 30784
rect 7607 30753 7619 30756
rect 7561 30747 7619 30753
rect 7377 30719 7435 30725
rect 7377 30685 7389 30719
rect 7423 30716 7435 30719
rect 7650 30716 7656 30728
rect 7423 30688 7656 30716
rect 7423 30685 7435 30688
rect 7377 30679 7435 30685
rect 7650 30676 7656 30688
rect 7708 30676 7714 30728
rect 9048 30580 9076 30756
rect 9122 30744 9128 30796
rect 9180 30784 9186 30796
rect 10781 30787 10839 30793
rect 10781 30784 10793 30787
rect 9180 30756 10793 30784
rect 9180 30744 9186 30756
rect 10781 30753 10793 30756
rect 10827 30784 10839 30787
rect 13464 30784 13492 30824
rect 10827 30756 13492 30784
rect 13541 30787 13599 30793
rect 10827 30753 10839 30756
rect 10781 30747 10839 30753
rect 13541 30753 13553 30787
rect 13587 30753 13599 30787
rect 13541 30747 13599 30753
rect 10318 30608 10324 30660
rect 10376 30648 10382 30660
rect 13556 30648 13584 30747
rect 14292 30728 14320 30824
rect 17034 30812 17040 30864
rect 17092 30852 17098 30864
rect 24857 30855 24915 30861
rect 17092 30824 17632 30852
rect 17092 30812 17098 30824
rect 17310 30744 17316 30796
rect 17368 30784 17374 30796
rect 17604 30793 17632 30824
rect 24857 30821 24869 30855
rect 24903 30852 24915 30855
rect 25958 30852 25964 30864
rect 24903 30824 25964 30852
rect 24903 30821 24915 30824
rect 24857 30815 24915 30821
rect 25958 30812 25964 30824
rect 26016 30812 26022 30864
rect 17497 30787 17555 30793
rect 17497 30784 17509 30787
rect 17368 30756 17509 30784
rect 17368 30744 17374 30756
rect 17497 30753 17509 30756
rect 17543 30753 17555 30787
rect 17497 30747 17555 30753
rect 17589 30787 17647 30793
rect 17589 30753 17601 30787
rect 17635 30753 17647 30787
rect 17589 30747 17647 30753
rect 22281 30787 22339 30793
rect 22281 30753 22293 30787
rect 22327 30784 22339 30787
rect 22646 30784 22652 30796
rect 22327 30756 22652 30784
rect 22327 30753 22339 30756
rect 22281 30747 22339 30753
rect 22646 30744 22652 30756
rect 22704 30744 22710 30796
rect 24210 30784 24216 30796
rect 23676 30756 24216 30784
rect 14274 30676 14280 30728
rect 14332 30676 14338 30728
rect 17402 30676 17408 30728
rect 17460 30676 17466 30728
rect 23676 30702 23704 30756
rect 24210 30744 24216 30756
rect 24268 30784 24274 30796
rect 24486 30784 24492 30796
rect 24268 30756 24492 30784
rect 24268 30744 24274 30756
rect 24486 30744 24492 30756
rect 24544 30744 24550 30796
rect 10376 30620 11546 30648
rect 12360 30620 13584 30648
rect 10376 30608 10382 30620
rect 9398 30580 9404 30592
rect 9048 30552 9404 30580
rect 9398 30540 9404 30552
rect 9456 30580 9462 30592
rect 12360 30580 12388 30620
rect 14458 30608 14464 30660
rect 14516 30648 14522 30660
rect 14553 30651 14611 30657
rect 14553 30648 14565 30651
rect 14516 30620 14565 30648
rect 14516 30608 14522 30620
rect 14553 30617 14565 30620
rect 14599 30617 14611 30651
rect 14553 30611 14611 30617
rect 15194 30608 15200 30660
rect 15252 30608 15258 30660
rect 22462 30608 22468 30660
rect 22520 30648 22526 30660
rect 22557 30651 22615 30657
rect 22557 30648 22569 30651
rect 22520 30620 22569 30648
rect 22520 30608 22526 30620
rect 22557 30617 22569 30620
rect 22603 30617 22615 30651
rect 22557 30611 22615 30617
rect 24486 30608 24492 30660
rect 24544 30648 24550 30660
rect 24673 30651 24731 30657
rect 24673 30648 24685 30651
rect 24544 30620 24685 30648
rect 24544 30608 24550 30620
rect 24673 30617 24685 30620
rect 24719 30617 24731 30651
rect 24673 30611 24731 30617
rect 9456 30552 12388 30580
rect 9456 30540 9462 30552
rect 12526 30540 12532 30592
rect 12584 30540 12590 30592
rect 12618 30540 12624 30592
rect 12676 30580 12682 30592
rect 13354 30580 13360 30592
rect 12676 30552 13360 30580
rect 12676 30540 12682 30552
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 13449 30583 13507 30589
rect 13449 30549 13461 30583
rect 13495 30580 13507 30583
rect 14182 30580 14188 30592
rect 13495 30552 14188 30580
rect 13495 30549 13507 30552
rect 13449 30543 13507 30549
rect 14182 30540 14188 30552
rect 14240 30540 14246 30592
rect 15930 30540 15936 30592
rect 15988 30580 15994 30592
rect 16025 30583 16083 30589
rect 16025 30580 16037 30583
rect 15988 30552 16037 30580
rect 15988 30540 15994 30552
rect 16025 30549 16037 30552
rect 16071 30580 16083 30583
rect 16206 30580 16212 30592
rect 16071 30552 16212 30580
rect 16071 30549 16083 30552
rect 16025 30543 16083 30549
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 16666 30540 16672 30592
rect 16724 30580 16730 30592
rect 17037 30583 17095 30589
rect 17037 30580 17049 30583
rect 16724 30552 17049 30580
rect 16724 30540 16730 30552
rect 17037 30549 17049 30552
rect 17083 30549 17095 30583
rect 17037 30543 17095 30549
rect 24026 30540 24032 30592
rect 24084 30540 24090 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 9030 30376 9036 30388
rect 8312 30348 9036 30376
rect 8312 30308 8340 30348
rect 9030 30336 9036 30348
rect 9088 30336 9094 30388
rect 13354 30336 13360 30388
rect 13412 30376 13418 30388
rect 16942 30376 16948 30388
rect 13412 30348 16948 30376
rect 13412 30336 13418 30348
rect 16942 30336 16948 30348
rect 17000 30336 17006 30388
rect 25038 30376 25044 30388
rect 20824 30348 25044 30376
rect 20824 30320 20852 30348
rect 25038 30336 25044 30348
rect 25096 30336 25102 30388
rect 10318 30308 10324 30320
rect 7760 30280 8340 30308
rect 9246 30280 10324 30308
rect 7760 30249 7788 30280
rect 10318 30268 10324 30280
rect 10376 30268 10382 30320
rect 13081 30311 13139 30317
rect 13081 30277 13093 30311
rect 13127 30308 13139 30311
rect 15010 30308 15016 30320
rect 13127 30280 15016 30308
rect 13127 30277 13139 30280
rect 13081 30271 13139 30277
rect 15010 30268 15016 30280
rect 15068 30268 15074 30320
rect 15197 30311 15255 30317
rect 15197 30277 15209 30311
rect 15243 30308 15255 30311
rect 18506 30308 18512 30320
rect 15243 30280 18512 30308
rect 15243 30277 15255 30280
rect 15197 30271 15255 30277
rect 18506 30268 18512 30280
rect 18564 30268 18570 30320
rect 18598 30268 18604 30320
rect 18656 30308 18662 30320
rect 18966 30308 18972 30320
rect 18656 30280 18972 30308
rect 18656 30268 18662 30280
rect 18966 30268 18972 30280
rect 19024 30268 19030 30320
rect 19886 30268 19892 30320
rect 19944 30308 19950 30320
rect 20438 30308 20444 30320
rect 19944 30280 20444 30308
rect 19944 30268 19950 30280
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 20806 30268 20812 30320
rect 20864 30268 20870 30320
rect 20901 30311 20959 30317
rect 20901 30277 20913 30311
rect 20947 30308 20959 30311
rect 21358 30308 21364 30320
rect 20947 30280 21364 30308
rect 20947 30277 20959 30280
rect 20901 30271 20959 30277
rect 21358 30268 21364 30280
rect 21416 30268 21422 30320
rect 22278 30268 22284 30320
rect 22336 30308 22342 30320
rect 22373 30311 22431 30317
rect 22373 30308 22385 30311
rect 22336 30280 22385 30308
rect 22336 30268 22342 30280
rect 22373 30277 22385 30280
rect 22419 30277 22431 30311
rect 22373 30271 22431 30277
rect 24210 30268 24216 30320
rect 24268 30268 24274 30320
rect 7745 30243 7803 30249
rect 7745 30209 7757 30243
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 12986 30200 12992 30252
rect 13044 30200 13050 30252
rect 14366 30200 14372 30252
rect 14424 30240 14430 30252
rect 17221 30243 17279 30249
rect 17221 30240 17233 30243
rect 14424 30212 17233 30240
rect 14424 30200 14430 30212
rect 17221 30209 17233 30212
rect 17267 30209 17279 30243
rect 17221 30203 17279 30209
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30240 17371 30243
rect 19150 30240 19156 30252
rect 17359 30212 19156 30240
rect 17359 30209 17371 30212
rect 17313 30203 17371 30209
rect 19150 30200 19156 30212
rect 19208 30200 19214 30252
rect 19613 30243 19671 30249
rect 19613 30209 19625 30243
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 19705 30243 19763 30249
rect 19705 30209 19717 30243
rect 19751 30240 19763 30243
rect 20162 30240 20168 30252
rect 19751 30212 20168 30240
rect 19751 30209 19763 30212
rect 19705 30203 19763 30209
rect 8018 30132 8024 30184
rect 8076 30132 8082 30184
rect 8386 30132 8392 30184
rect 8444 30172 8450 30184
rect 9493 30175 9551 30181
rect 9493 30172 9505 30175
rect 8444 30144 9505 30172
rect 8444 30132 8450 30144
rect 9493 30141 9505 30144
rect 9539 30141 9551 30175
rect 9493 30135 9551 30141
rect 9674 30132 9680 30184
rect 9732 30172 9738 30184
rect 13265 30175 13323 30181
rect 9732 30144 13032 30172
rect 9732 30132 9738 30144
rect 10410 30064 10416 30116
rect 10468 30104 10474 30116
rect 12621 30107 12679 30113
rect 12621 30104 12633 30107
rect 10468 30076 12633 30104
rect 10468 30064 10474 30076
rect 12621 30073 12633 30076
rect 12667 30073 12679 30107
rect 13004 30104 13032 30144
rect 13265 30141 13277 30175
rect 13311 30172 13323 30175
rect 14642 30172 14648 30184
rect 13311 30144 14648 30172
rect 13311 30141 13323 30144
rect 13265 30135 13323 30141
rect 13280 30104 13308 30135
rect 14642 30132 14648 30144
rect 14700 30132 14706 30184
rect 15286 30132 15292 30184
rect 15344 30132 15350 30184
rect 15381 30175 15439 30181
rect 15381 30141 15393 30175
rect 15427 30141 15439 30175
rect 15381 30135 15439 30141
rect 13004 30076 13308 30104
rect 12621 30067 12679 30073
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 15396 30104 15424 30135
rect 16942 30132 16948 30184
rect 17000 30172 17006 30184
rect 17405 30175 17463 30181
rect 17405 30172 17417 30175
rect 17000 30144 17417 30172
rect 17000 30132 17006 30144
rect 17405 30141 17417 30144
rect 17451 30172 17463 30175
rect 17586 30172 17592 30184
rect 17451 30144 17592 30172
rect 17451 30141 17463 30144
rect 17405 30135 17463 30141
rect 17586 30132 17592 30144
rect 17644 30132 17650 30184
rect 19628 30172 19656 30203
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 21726 30200 21732 30252
rect 21784 30240 21790 30252
rect 21784 30212 22094 30240
rect 21784 30200 21790 30212
rect 18432 30144 19656 30172
rect 19889 30175 19947 30181
rect 14056 30076 15424 30104
rect 16316 30076 17448 30104
rect 14056 30064 14062 30076
rect 3602 29996 3608 30048
rect 3660 30036 3666 30048
rect 8478 30036 8484 30048
rect 3660 30008 8484 30036
rect 3660 29996 3666 30008
rect 8478 29996 8484 30008
rect 8536 30036 8542 30048
rect 9398 30036 9404 30048
rect 8536 30008 9404 30036
rect 8536 29996 8542 30008
rect 9398 29996 9404 30008
rect 9456 29996 9462 30048
rect 10962 29996 10968 30048
rect 11020 30036 11026 30048
rect 11885 30039 11943 30045
rect 11885 30036 11897 30039
rect 11020 30008 11897 30036
rect 11020 29996 11026 30008
rect 11885 30005 11897 30008
rect 11931 30005 11943 30039
rect 11885 29999 11943 30005
rect 13538 29996 13544 30048
rect 13596 30036 13602 30048
rect 14829 30039 14887 30045
rect 14829 30036 14841 30039
rect 13596 30008 14841 30036
rect 13596 29996 13602 30008
rect 14829 30005 14841 30008
rect 14875 30005 14887 30039
rect 14829 29999 14887 30005
rect 14918 29996 14924 30048
rect 14976 30036 14982 30048
rect 16316 30036 16344 30076
rect 14976 30008 16344 30036
rect 16853 30039 16911 30045
rect 14976 29996 14982 30008
rect 16853 30005 16865 30039
rect 16899 30036 16911 30039
rect 17310 30036 17316 30048
rect 16899 30008 17316 30036
rect 16899 30005 16911 30008
rect 16853 29999 16911 30005
rect 17310 29996 17316 30008
rect 17368 29996 17374 30048
rect 17420 30036 17448 30076
rect 18432 30036 18460 30144
rect 19889 30141 19901 30175
rect 19935 30172 19947 30175
rect 20254 30172 20260 30184
rect 19935 30144 20260 30172
rect 19935 30141 19947 30144
rect 19889 30135 19947 30141
rect 20254 30132 20260 30144
rect 20312 30132 20318 30184
rect 20993 30175 21051 30181
rect 20993 30172 21005 30175
rect 20364 30144 21005 30172
rect 18506 30064 18512 30116
rect 18564 30104 18570 30116
rect 19245 30107 19303 30113
rect 18564 30076 18828 30104
rect 18564 30064 18570 30076
rect 18693 30039 18751 30045
rect 18693 30036 18705 30039
rect 17420 30008 18705 30036
rect 18693 30005 18705 30008
rect 18739 30005 18751 30039
rect 18800 30036 18828 30076
rect 19245 30073 19257 30107
rect 19291 30104 19303 30107
rect 19426 30104 19432 30116
rect 19291 30076 19432 30104
rect 19291 30073 19303 30076
rect 19245 30067 19303 30073
rect 19426 30064 19432 30076
rect 19484 30064 19490 30116
rect 20364 30036 20392 30144
rect 20993 30141 21005 30144
rect 21039 30141 21051 30175
rect 22066 30172 22094 30212
rect 22646 30200 22652 30252
rect 22704 30240 22710 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22704 30212 23397 30240
rect 22704 30200 22710 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 22465 30175 22523 30181
rect 22465 30172 22477 30175
rect 22066 30144 22477 30172
rect 20993 30135 21051 30141
rect 22465 30141 22477 30144
rect 22511 30141 22523 30175
rect 22465 30135 22523 30141
rect 22557 30175 22615 30181
rect 22557 30141 22569 30175
rect 22603 30172 22615 30175
rect 23661 30175 23719 30181
rect 23661 30172 23673 30175
rect 22603 30144 23673 30172
rect 22603 30141 22615 30144
rect 22557 30135 22615 30141
rect 23661 30141 23673 30144
rect 23707 30172 23719 30175
rect 24026 30172 24032 30184
rect 23707 30144 24032 30172
rect 23707 30141 23719 30144
rect 23661 30135 23719 30141
rect 22572 30104 22600 30135
rect 24026 30132 24032 30144
rect 24084 30132 24090 30184
rect 22646 30104 22652 30116
rect 22572 30076 22652 30104
rect 22646 30064 22652 30076
rect 22704 30064 22710 30116
rect 18800 30008 20392 30036
rect 18693 29999 18751 30005
rect 20438 29996 20444 30048
rect 20496 29996 20502 30048
rect 22005 30039 22063 30045
rect 22005 30005 22017 30039
rect 22051 30036 22063 30039
rect 23474 30036 23480 30048
rect 22051 30008 23480 30036
rect 22051 30005 22063 30008
rect 22005 29999 22063 30005
rect 23474 29996 23480 30008
rect 23532 29996 23538 30048
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 25133 30039 25191 30045
rect 25133 30036 25145 30039
rect 23808 30008 25145 30036
rect 23808 29996 23814 30008
rect 25133 30005 25145 30008
rect 25179 30005 25191 30039
rect 25133 29999 25191 30005
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 8938 29792 8944 29844
rect 8996 29832 9002 29844
rect 9125 29835 9183 29841
rect 9125 29832 9137 29835
rect 8996 29804 9137 29832
rect 8996 29792 9002 29804
rect 9125 29801 9137 29804
rect 9171 29801 9183 29835
rect 12618 29832 12624 29844
rect 9125 29795 9183 29801
rect 10060 29804 12624 29832
rect 7558 29724 7564 29776
rect 7616 29764 7622 29776
rect 9674 29764 9680 29776
rect 7616 29736 9680 29764
rect 7616 29724 7622 29736
rect 9674 29724 9680 29736
rect 9732 29724 9738 29776
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1360 29668 2053 29696
rect 1360 29656 1366 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 8018 29656 8024 29708
rect 8076 29696 8082 29708
rect 9766 29696 9772 29708
rect 8076 29668 9772 29696
rect 8076 29656 8082 29668
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 1762 29588 1768 29640
rect 1820 29588 1826 29640
rect 1854 29588 1860 29640
rect 1912 29628 1918 29640
rect 3973 29631 4031 29637
rect 3973 29628 3985 29631
rect 1912 29600 3985 29628
rect 1912 29588 1918 29600
rect 3973 29597 3985 29600
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 9398 29588 9404 29640
rect 9456 29628 9462 29640
rect 9493 29631 9551 29637
rect 9493 29628 9505 29631
rect 9456 29600 9505 29628
rect 9456 29588 9462 29600
rect 9493 29597 9505 29600
rect 9539 29597 9551 29631
rect 10060 29628 10088 29804
rect 12618 29792 12624 29804
rect 12676 29832 12682 29844
rect 13354 29832 13360 29844
rect 12676 29804 13360 29832
rect 12676 29792 12682 29804
rect 13354 29792 13360 29804
rect 13412 29792 13418 29844
rect 14090 29792 14096 29844
rect 14148 29832 14154 29844
rect 14918 29832 14924 29844
rect 14148 29804 14924 29832
rect 14148 29792 14154 29804
rect 14918 29792 14924 29804
rect 14976 29792 14982 29844
rect 17129 29835 17187 29841
rect 17129 29801 17141 29835
rect 17175 29832 17187 29835
rect 19242 29832 19248 29844
rect 17175 29804 19248 29832
rect 17175 29801 17187 29804
rect 17129 29795 17187 29801
rect 19242 29792 19248 29804
rect 19300 29792 19306 29844
rect 22462 29832 22468 29844
rect 22066 29804 22468 29832
rect 10410 29724 10416 29776
rect 10468 29764 10474 29776
rect 11793 29767 11851 29773
rect 11793 29764 11805 29767
rect 10468 29736 11805 29764
rect 10468 29724 10474 29736
rect 11793 29733 11805 29736
rect 11839 29733 11851 29767
rect 11793 29727 11851 29733
rect 12158 29724 12164 29776
rect 12216 29764 12222 29776
rect 18049 29767 18107 29773
rect 18049 29764 18061 29767
rect 12216 29736 18061 29764
rect 12216 29724 12222 29736
rect 18049 29733 18061 29736
rect 18095 29733 18107 29767
rect 19610 29764 19616 29776
rect 18049 29727 18107 29733
rect 18156 29736 19616 29764
rect 10134 29656 10140 29708
rect 10192 29696 10198 29708
rect 10594 29696 10600 29708
rect 10192 29668 10600 29696
rect 10192 29656 10198 29668
rect 10594 29656 10600 29668
rect 10652 29696 10658 29708
rect 11057 29699 11115 29705
rect 11057 29696 11069 29699
rect 10652 29668 11069 29696
rect 10652 29656 10658 29668
rect 11057 29665 11069 29668
rect 11103 29665 11115 29699
rect 11057 29659 11115 29665
rect 11238 29656 11244 29708
rect 11296 29656 11302 29708
rect 12253 29699 12311 29705
rect 12253 29696 12265 29699
rect 12176 29668 12265 29696
rect 12176 29640 12204 29668
rect 12253 29665 12265 29668
rect 12299 29665 12311 29699
rect 12253 29659 12311 29665
rect 12345 29699 12403 29705
rect 12345 29665 12357 29699
rect 12391 29696 12403 29699
rect 12434 29696 12440 29708
rect 12391 29668 12440 29696
rect 12391 29665 12403 29668
rect 12345 29659 12403 29665
rect 12434 29656 12440 29668
rect 12492 29656 12498 29708
rect 13446 29656 13452 29708
rect 13504 29656 13510 29708
rect 13541 29699 13599 29705
rect 13541 29665 13553 29699
rect 13587 29665 13599 29699
rect 13541 29659 13599 29665
rect 17773 29699 17831 29705
rect 17773 29665 17785 29699
rect 17819 29696 17831 29699
rect 18156 29696 18184 29736
rect 19610 29724 19616 29736
rect 19668 29764 19674 29776
rect 20714 29764 20720 29776
rect 19668 29736 20720 29764
rect 19668 29724 19674 29736
rect 20714 29724 20720 29736
rect 20772 29724 20778 29776
rect 21266 29724 21272 29776
rect 21324 29764 21330 29776
rect 21913 29767 21971 29773
rect 21324 29736 21864 29764
rect 21324 29724 21330 29736
rect 17819 29668 18184 29696
rect 18601 29699 18659 29705
rect 17819 29665 17831 29668
rect 17773 29659 17831 29665
rect 18601 29665 18613 29699
rect 18647 29665 18659 29699
rect 18601 29659 18659 29665
rect 9493 29591 9551 29597
rect 9600 29600 10088 29628
rect 3510 29520 3516 29572
rect 3568 29560 3574 29572
rect 4157 29563 4215 29569
rect 4157 29560 4169 29563
rect 3568 29532 4169 29560
rect 3568 29520 3574 29532
rect 4157 29529 4169 29532
rect 4203 29529 4215 29563
rect 4157 29523 4215 29529
rect 5813 29563 5871 29569
rect 5813 29529 5825 29563
rect 5859 29560 5871 29563
rect 5994 29560 6000 29572
rect 5859 29532 6000 29560
rect 5859 29529 5871 29532
rect 5813 29523 5871 29529
rect 5994 29520 6000 29532
rect 6052 29520 6058 29572
rect 8846 29520 8852 29572
rect 8904 29560 8910 29572
rect 9600 29569 9628 29600
rect 10962 29588 10968 29640
rect 11020 29588 11026 29640
rect 12158 29588 12164 29640
rect 12216 29588 12222 29640
rect 13357 29631 13415 29637
rect 13357 29628 13369 29631
rect 12268 29600 13369 29628
rect 9585 29563 9643 29569
rect 9585 29560 9597 29563
rect 8904 29532 9597 29560
rect 8904 29520 8910 29532
rect 9585 29529 9597 29532
rect 9631 29529 9643 29563
rect 12268 29560 12296 29600
rect 13357 29597 13369 29600
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 9585 29523 9643 29529
rect 10612 29532 12296 29560
rect 10612 29501 10640 29532
rect 12526 29520 12532 29572
rect 12584 29560 12590 29572
rect 13556 29560 13584 29659
rect 14826 29588 14832 29640
rect 14884 29628 14890 29640
rect 18616 29628 18644 29659
rect 19334 29656 19340 29708
rect 19392 29696 19398 29708
rect 19889 29699 19947 29705
rect 19889 29696 19901 29699
rect 19392 29668 19901 29696
rect 19392 29656 19398 29668
rect 19889 29665 19901 29668
rect 19935 29665 19947 29699
rect 19889 29659 19947 29665
rect 19981 29699 20039 29705
rect 19981 29665 19993 29699
rect 20027 29665 20039 29699
rect 19981 29659 20039 29665
rect 14884 29600 18644 29628
rect 14884 29588 14890 29600
rect 18690 29588 18696 29640
rect 18748 29628 18754 29640
rect 19996 29628 20024 29659
rect 21174 29656 21180 29708
rect 21232 29656 21238 29708
rect 21361 29699 21419 29705
rect 21361 29665 21373 29699
rect 21407 29696 21419 29699
rect 21726 29696 21732 29708
rect 21407 29668 21732 29696
rect 21407 29665 21419 29668
rect 21361 29659 21419 29665
rect 21726 29656 21732 29668
rect 21784 29656 21790 29708
rect 21836 29696 21864 29736
rect 21913 29733 21925 29767
rect 21959 29764 21971 29767
rect 22066 29764 22094 29804
rect 22462 29792 22468 29804
rect 22520 29792 22526 29844
rect 25130 29792 25136 29844
rect 25188 29792 25194 29844
rect 21959 29736 22094 29764
rect 23109 29767 23167 29773
rect 21959 29733 21971 29736
rect 21913 29727 21971 29733
rect 23109 29733 23121 29767
rect 23155 29764 23167 29767
rect 24026 29764 24032 29776
rect 23155 29736 24032 29764
rect 23155 29733 23167 29736
rect 23109 29727 23167 29733
rect 24026 29724 24032 29736
rect 24084 29724 24090 29776
rect 22465 29699 22523 29705
rect 22465 29696 22477 29699
rect 21836 29668 22477 29696
rect 22465 29665 22477 29668
rect 22511 29665 22523 29699
rect 22465 29659 22523 29665
rect 23474 29656 23480 29708
rect 23532 29696 23538 29708
rect 23569 29699 23627 29705
rect 23569 29696 23581 29699
rect 23532 29668 23581 29696
rect 23532 29656 23538 29668
rect 23569 29665 23581 29668
rect 23615 29665 23627 29699
rect 23569 29659 23627 29665
rect 23750 29656 23756 29708
rect 23808 29656 23814 29708
rect 18748 29600 20024 29628
rect 21085 29631 21143 29637
rect 18748 29588 18754 29600
rect 21085 29597 21097 29631
rect 21131 29628 21143 29631
rect 22186 29628 22192 29640
rect 21131 29600 22192 29628
rect 21131 29597 21143 29600
rect 21085 29591 21143 29597
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 22370 29588 22376 29640
rect 22428 29588 22434 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 18322 29560 18328 29572
rect 12584 29532 13584 29560
rect 17420 29532 18328 29560
rect 12584 29520 12590 29532
rect 10597 29495 10655 29501
rect 10597 29461 10609 29495
rect 10643 29461 10655 29495
rect 10597 29455 10655 29461
rect 12161 29495 12219 29501
rect 12161 29461 12173 29495
rect 12207 29492 12219 29495
rect 12894 29492 12900 29504
rect 12207 29464 12900 29492
rect 12207 29461 12219 29464
rect 12161 29455 12219 29461
rect 12894 29452 12900 29464
rect 12952 29452 12958 29504
rect 12989 29495 13047 29501
rect 12989 29461 13001 29495
rect 13035 29492 13047 29495
rect 17420 29492 17448 29532
rect 18322 29520 18328 29532
rect 18380 29520 18386 29572
rect 18509 29563 18567 29569
rect 18509 29529 18521 29563
rect 18555 29560 18567 29563
rect 22281 29563 22339 29569
rect 22281 29560 22293 29563
rect 18555 29532 22293 29560
rect 18555 29529 18567 29532
rect 18509 29523 18567 29529
rect 22281 29529 22293 29532
rect 22327 29560 22339 29563
rect 23566 29560 23572 29572
rect 22327 29532 23572 29560
rect 22327 29529 22339 29532
rect 22281 29523 22339 29529
rect 23566 29520 23572 29532
rect 23624 29520 23630 29572
rect 13035 29464 17448 29492
rect 13035 29461 13047 29464
rect 12989 29455 13047 29461
rect 17494 29452 17500 29504
rect 17552 29452 17558 29504
rect 17586 29452 17592 29504
rect 17644 29452 17650 29504
rect 18417 29495 18475 29501
rect 18417 29461 18429 29495
rect 18463 29492 18475 29495
rect 18966 29492 18972 29504
rect 18463 29464 18972 29492
rect 18463 29461 18475 29464
rect 18417 29455 18475 29461
rect 18966 29452 18972 29464
rect 19024 29452 19030 29504
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19392 29464 19441 29492
rect 19392 29452 19398 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19797 29495 19855 29501
rect 19797 29461 19809 29495
rect 19843 29492 19855 29495
rect 19978 29492 19984 29504
rect 19843 29464 19984 29492
rect 19843 29461 19855 29464
rect 19797 29455 19855 29461
rect 19978 29452 19984 29464
rect 20036 29452 20042 29504
rect 20717 29495 20775 29501
rect 20717 29461 20729 29495
rect 20763 29492 20775 29495
rect 20990 29492 20996 29504
rect 20763 29464 20996 29492
rect 20763 29461 20775 29464
rect 20717 29455 20775 29461
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 23290 29452 23296 29504
rect 23348 29492 23354 29504
rect 23477 29495 23535 29501
rect 23477 29492 23489 29495
rect 23348 29464 23489 29492
rect 23348 29452 23354 29464
rect 23477 29461 23489 29464
rect 23523 29461 23535 29495
rect 23477 29455 23535 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8202 29248 8208 29300
rect 8260 29288 8266 29300
rect 9861 29291 9919 29297
rect 9861 29288 9873 29291
rect 8260 29260 9873 29288
rect 8260 29248 8266 29260
rect 9861 29257 9873 29260
rect 9907 29288 9919 29291
rect 12434 29288 12440 29300
rect 9907 29260 12440 29288
rect 9907 29257 9919 29260
rect 9861 29251 9919 29257
rect 12434 29248 12440 29260
rect 12492 29248 12498 29300
rect 13354 29248 13360 29300
rect 13412 29288 13418 29300
rect 13722 29288 13728 29300
rect 13412 29260 13728 29288
rect 13412 29248 13418 29260
rect 13722 29248 13728 29260
rect 13780 29288 13786 29300
rect 17494 29288 17500 29300
rect 13780 29260 17500 29288
rect 13780 29248 13786 29260
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 17604 29260 19472 29288
rect 8662 29220 8668 29232
rect 8128 29192 8668 29220
rect 8128 29161 8156 29192
rect 8662 29180 8668 29192
rect 8720 29180 8726 29232
rect 10318 29220 10324 29232
rect 9614 29192 10324 29220
rect 10318 29180 10324 29192
rect 10376 29180 10382 29232
rect 11146 29180 11152 29232
rect 11204 29220 11210 29232
rect 12253 29223 12311 29229
rect 12253 29220 12265 29223
rect 11204 29192 12265 29220
rect 11204 29180 11210 29192
rect 12253 29189 12265 29192
rect 12299 29220 12311 29223
rect 14366 29220 14372 29232
rect 12299 29192 14372 29220
rect 12299 29189 12311 29192
rect 12253 29183 12311 29189
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 17126 29220 17132 29232
rect 14476 29192 17132 29220
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29121 8171 29155
rect 8113 29115 8171 29121
rect 12161 29155 12219 29161
rect 12161 29121 12173 29155
rect 12207 29152 12219 29155
rect 14476 29152 14504 29192
rect 17126 29180 17132 29192
rect 17184 29180 17190 29232
rect 12207 29124 14504 29152
rect 12207 29121 12219 29124
rect 12161 29115 12219 29121
rect 14550 29112 14556 29164
rect 14608 29112 14614 29164
rect 17604 29152 17632 29260
rect 19058 29180 19064 29232
rect 19116 29180 19122 29232
rect 19444 29220 19472 29260
rect 19518 29248 19524 29300
rect 19576 29288 19582 29300
rect 21082 29288 21088 29300
rect 19576 29260 21088 29288
rect 19576 29248 19582 29260
rect 21082 29248 21088 29260
rect 21140 29248 21146 29300
rect 20622 29220 20628 29232
rect 19444 29192 20628 29220
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24673 29223 24731 29229
rect 24673 29220 24685 29223
rect 24636 29192 24685 29220
rect 24636 29180 24642 29192
rect 24673 29189 24685 29192
rect 24719 29189 24731 29223
rect 24673 29183 24731 29189
rect 14936 29124 17632 29152
rect 17773 29155 17831 29161
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 12345 29087 12403 29093
rect 9732 29056 11928 29084
rect 9732 29044 9738 29056
rect 9784 28988 9996 29016
rect 8376 28951 8434 28957
rect 8376 28917 8388 28951
rect 8422 28948 8434 28951
rect 9784 28948 9812 28988
rect 8422 28920 9812 28948
rect 9968 28948 9996 28988
rect 10226 28976 10232 29028
rect 10284 29016 10290 29028
rect 11793 29019 11851 29025
rect 11793 29016 11805 29019
rect 10284 28988 11805 29016
rect 10284 28976 10290 28988
rect 11793 28985 11805 28988
rect 11839 28985 11851 29019
rect 11900 29016 11928 29056
rect 12345 29053 12357 29087
rect 12391 29053 12403 29087
rect 12345 29047 12403 29053
rect 12360 29016 12388 29047
rect 14936 29028 14964 29124
rect 17773 29121 17785 29155
rect 17819 29121 17831 29155
rect 17773 29115 17831 29121
rect 11900 28988 12388 29016
rect 11793 28979 11851 28985
rect 12434 28976 12440 29028
rect 12492 29016 12498 29028
rect 12618 29016 12624 29028
rect 12492 28988 12624 29016
rect 12492 28976 12498 28988
rect 12618 28976 12624 28988
rect 12676 28976 12682 29028
rect 12894 28976 12900 29028
rect 12952 29016 12958 29028
rect 14918 29016 14924 29028
rect 12952 28988 14924 29016
rect 12952 28976 12958 28988
rect 14918 28976 14924 28988
rect 14976 28976 14982 29028
rect 15838 28976 15844 29028
rect 15896 29016 15902 29028
rect 16022 29016 16028 29028
rect 15896 28988 16028 29016
rect 15896 28976 15902 28988
rect 16022 28976 16028 28988
rect 16080 28976 16086 29028
rect 16758 28976 16764 29028
rect 16816 29016 16822 29028
rect 17788 29016 17816 29115
rect 24118 29112 24124 29164
rect 24176 29112 24182 29164
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 19521 29087 19579 29093
rect 19521 29084 19533 29087
rect 18196 29056 19533 29084
rect 18196 29044 18202 29056
rect 19521 29053 19533 29056
rect 19567 29053 19579 29087
rect 19521 29047 19579 29053
rect 16816 28988 17816 29016
rect 16816 28976 16822 28988
rect 19058 28976 19064 29028
rect 19116 29016 19122 29028
rect 23937 29019 23995 29025
rect 23937 29016 23949 29019
rect 19116 28988 23949 29016
rect 19116 28976 19122 28988
rect 23937 28985 23949 28988
rect 23983 28985 23995 29019
rect 23937 28979 23995 28985
rect 24394 28976 24400 29028
rect 24452 29016 24458 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 24452 28988 24869 29016
rect 24452 28976 24458 28988
rect 24857 28985 24869 28988
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 11054 28948 11060 28960
rect 9968 28920 11060 28948
rect 8422 28917 8434 28920
rect 8376 28911 8434 28917
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 18036 28951 18094 28957
rect 18036 28917 18048 28951
rect 18082 28948 18094 28951
rect 18598 28948 18604 28960
rect 18082 28920 18604 28948
rect 18082 28917 18094 28920
rect 18036 28911 18094 28917
rect 18598 28908 18604 28920
rect 18656 28908 18662 28960
rect 22186 28908 22192 28960
rect 22244 28908 22250 28960
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 9125 28747 9183 28753
rect 9125 28713 9137 28747
rect 9171 28744 9183 28747
rect 9306 28744 9312 28756
rect 9171 28716 9312 28744
rect 9171 28713 9183 28716
rect 9125 28707 9183 28713
rect 9306 28704 9312 28716
rect 9364 28704 9370 28756
rect 9582 28704 9588 28756
rect 9640 28704 9646 28756
rect 15378 28704 15384 28756
rect 15436 28744 15442 28756
rect 16298 28744 16304 28756
rect 15436 28716 16304 28744
rect 15436 28704 15442 28716
rect 16298 28704 16304 28716
rect 16356 28704 16362 28756
rect 16482 28704 16488 28756
rect 16540 28744 16546 28756
rect 20073 28747 20131 28753
rect 20073 28744 20085 28747
rect 16540 28716 20085 28744
rect 16540 28704 16546 28716
rect 20073 28713 20085 28716
rect 20119 28744 20131 28747
rect 20806 28744 20812 28756
rect 20119 28716 20812 28744
rect 20119 28713 20131 28716
rect 20073 28707 20131 28713
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 21821 28747 21879 28753
rect 21821 28713 21833 28747
rect 21867 28744 21879 28747
rect 23290 28744 23296 28756
rect 21867 28716 23296 28744
rect 21867 28713 21879 28716
rect 21821 28707 21879 28713
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 23934 28704 23940 28756
rect 23992 28744 23998 28756
rect 25133 28747 25191 28753
rect 25133 28744 25145 28747
rect 23992 28716 25145 28744
rect 23992 28704 23998 28716
rect 25133 28713 25145 28716
rect 25179 28713 25191 28747
rect 25133 28707 25191 28713
rect 9600 28676 9628 28704
rect 9600 28648 9720 28676
rect 3418 28568 3424 28620
rect 3476 28608 3482 28620
rect 3973 28611 4031 28617
rect 3973 28608 3985 28611
rect 3476 28580 3985 28608
rect 3476 28568 3482 28580
rect 3973 28577 3985 28580
rect 4019 28577 4031 28611
rect 3973 28571 4031 28577
rect 6549 28611 6607 28617
rect 6549 28577 6561 28611
rect 6595 28608 6607 28611
rect 6914 28608 6920 28620
rect 6595 28580 6920 28608
rect 6595 28577 6607 28580
rect 6549 28571 6607 28577
rect 6914 28568 6920 28580
rect 6972 28608 6978 28620
rect 8202 28608 8208 28620
rect 6972 28580 8208 28608
rect 6972 28568 6978 28580
rect 8202 28568 8208 28580
rect 8260 28568 8266 28620
rect 8570 28568 8576 28620
rect 8628 28608 8634 28620
rect 9692 28617 9720 28648
rect 16390 28636 16396 28688
rect 16448 28676 16454 28688
rect 16448 28648 22324 28676
rect 16448 28636 16454 28648
rect 9585 28611 9643 28617
rect 9585 28608 9597 28611
rect 8628 28580 9597 28608
rect 8628 28568 8634 28580
rect 9585 28577 9597 28580
rect 9631 28577 9643 28611
rect 9585 28571 9643 28577
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 11517 28611 11575 28617
rect 11517 28577 11529 28611
rect 11563 28608 11575 28611
rect 12526 28608 12532 28620
rect 11563 28580 12532 28608
rect 11563 28577 11575 28580
rect 11517 28571 11575 28577
rect 12526 28568 12532 28580
rect 12584 28568 12590 28620
rect 14274 28568 14280 28620
rect 14332 28608 14338 28620
rect 14553 28611 14611 28617
rect 14553 28608 14565 28611
rect 14332 28580 14565 28608
rect 14332 28568 14338 28580
rect 14553 28577 14565 28580
rect 14599 28577 14611 28611
rect 14553 28571 14611 28577
rect 14829 28611 14887 28617
rect 14829 28577 14841 28611
rect 14875 28608 14887 28611
rect 17497 28611 17555 28617
rect 17497 28608 17509 28611
rect 14875 28580 17509 28608
rect 14875 28577 14887 28580
rect 14829 28571 14887 28577
rect 17497 28577 17509 28580
rect 17543 28608 17555 28611
rect 17862 28608 17868 28620
rect 17543 28580 17868 28608
rect 17543 28577 17555 28580
rect 17497 28571 17555 28577
rect 17862 28568 17868 28580
rect 17920 28568 17926 28620
rect 20714 28568 20720 28620
rect 20772 28608 20778 28620
rect 20898 28608 20904 28620
rect 20772 28580 20904 28608
rect 20772 28568 20778 28580
rect 20898 28568 20904 28580
rect 20956 28608 20962 28620
rect 21085 28611 21143 28617
rect 21085 28608 21097 28611
rect 20956 28580 21097 28608
rect 20956 28568 20962 28580
rect 21085 28577 21097 28580
rect 21131 28577 21143 28611
rect 21085 28571 21143 28577
rect 21174 28568 21180 28620
rect 21232 28568 21238 28620
rect 22296 28617 22324 28648
rect 22281 28611 22339 28617
rect 22281 28577 22293 28611
rect 22327 28577 22339 28611
rect 22281 28571 22339 28577
rect 22465 28611 22523 28617
rect 22465 28577 22477 28611
rect 22511 28608 22523 28611
rect 22646 28608 22652 28620
rect 22511 28580 22652 28608
rect 22511 28577 22523 28580
rect 22465 28571 22523 28577
rect 22646 28568 22652 28580
rect 22704 28568 22710 28620
rect 6270 28500 6276 28552
rect 6328 28500 6334 28552
rect 8662 28500 8668 28552
rect 8720 28540 8726 28552
rect 11238 28540 11244 28552
rect 8720 28512 11244 28540
rect 8720 28500 8726 28512
rect 11238 28500 11244 28512
rect 11296 28500 11302 28552
rect 12618 28500 12624 28552
rect 12676 28500 12682 28552
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28540 17371 28543
rect 18325 28543 18383 28549
rect 18325 28540 18337 28543
rect 17359 28512 18337 28540
rect 17359 28509 17371 28512
rect 17313 28503 17371 28509
rect 18325 28509 18337 28512
rect 18371 28509 18383 28543
rect 18325 28503 18383 28509
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20346 28540 20352 28552
rect 20036 28512 20352 28540
rect 20036 28500 20042 28512
rect 20346 28500 20352 28512
rect 20404 28540 20410 28552
rect 20404 28512 22094 28540
rect 20404 28500 20410 28512
rect 4157 28475 4215 28481
rect 4157 28472 4169 28475
rect 3988 28444 4169 28472
rect 3988 28416 4016 28444
rect 4157 28441 4169 28444
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 5810 28432 5816 28484
rect 5868 28432 5874 28484
rect 7282 28432 7288 28484
rect 7340 28432 7346 28484
rect 8754 28472 8760 28484
rect 7944 28444 8760 28472
rect 3970 28364 3976 28416
rect 4028 28364 4034 28416
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 7944 28404 7972 28444
rect 8754 28432 8760 28444
rect 8812 28472 8818 28484
rect 9493 28475 9551 28481
rect 9493 28472 9505 28475
rect 8812 28444 9505 28472
rect 8812 28432 8818 28444
rect 9493 28441 9505 28444
rect 9539 28441 9551 28475
rect 9493 28435 9551 28441
rect 15378 28432 15384 28484
rect 15436 28432 15442 28484
rect 22066 28472 22094 28512
rect 22186 28500 22192 28552
rect 22244 28500 22250 28552
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28540 24087 28543
rect 24854 28540 24860 28552
rect 24075 28512 24860 28540
rect 24075 28509 24087 28512
rect 24029 28503 24087 28509
rect 24854 28500 24860 28512
rect 24912 28500 24918 28552
rect 25314 28500 25320 28552
rect 25372 28500 25378 28552
rect 20640 28444 21956 28472
rect 22066 28444 23888 28472
rect 4120 28376 7972 28404
rect 8021 28407 8079 28413
rect 4120 28364 4126 28376
rect 8021 28373 8033 28407
rect 8067 28404 8079 28407
rect 8294 28404 8300 28416
rect 8067 28376 8300 28404
rect 8067 28373 8079 28376
rect 8021 28367 8079 28373
rect 8294 28364 8300 28376
rect 8352 28364 8358 28416
rect 12802 28364 12808 28416
rect 12860 28404 12866 28416
rect 12989 28407 13047 28413
rect 12989 28404 13001 28407
rect 12860 28376 13001 28404
rect 12860 28364 12866 28376
rect 12989 28373 13001 28376
rect 13035 28373 13047 28407
rect 12989 28367 13047 28373
rect 16942 28364 16948 28416
rect 17000 28364 17006 28416
rect 17402 28364 17408 28416
rect 17460 28364 17466 28416
rect 20640 28413 20668 28444
rect 20625 28407 20683 28413
rect 20625 28373 20637 28407
rect 20671 28373 20683 28407
rect 20625 28367 20683 28373
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20864 28376 21005 28404
rect 20864 28364 20870 28376
rect 20993 28373 21005 28376
rect 21039 28373 21051 28407
rect 21928 28404 21956 28444
rect 22646 28404 22652 28416
rect 21928 28376 22652 28404
rect 20993 28367 21051 28373
rect 22646 28364 22652 28376
rect 22704 28364 22710 28416
rect 23860 28413 23888 28444
rect 23845 28407 23903 28413
rect 23845 28373 23857 28407
rect 23891 28373 23903 28407
rect 23845 28367 23903 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 7834 28160 7840 28212
rect 7892 28200 7898 28212
rect 8297 28203 8355 28209
rect 8297 28200 8309 28203
rect 7892 28172 8309 28200
rect 7892 28160 7898 28172
rect 8297 28169 8309 28172
rect 8343 28200 8355 28203
rect 9674 28200 9680 28212
rect 8343 28172 9680 28200
rect 8343 28169 8355 28172
rect 8297 28163 8355 28169
rect 9674 28160 9680 28172
rect 9732 28160 9738 28212
rect 10318 28160 10324 28212
rect 10376 28200 10382 28212
rect 10965 28203 11023 28209
rect 10376 28172 10640 28200
rect 10376 28160 10382 28172
rect 7282 28092 7288 28144
rect 7340 28092 7346 28144
rect 8662 28024 8668 28076
rect 8720 28064 8726 28076
rect 9217 28067 9275 28073
rect 9217 28064 9229 28067
rect 8720 28036 9229 28064
rect 8720 28024 8726 28036
rect 9217 28033 9229 28036
rect 9263 28033 9275 28067
rect 10612 28064 10640 28172
rect 10965 28169 10977 28203
rect 11011 28200 11023 28203
rect 11054 28200 11060 28212
rect 11011 28172 11060 28200
rect 11011 28169 11023 28172
rect 10965 28163 11023 28169
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 12342 28160 12348 28212
rect 12400 28160 12406 28212
rect 17310 28160 17316 28212
rect 17368 28160 17374 28212
rect 17402 28160 17408 28212
rect 17460 28200 17466 28212
rect 18049 28203 18107 28209
rect 18049 28200 18061 28203
rect 17460 28172 18061 28200
rect 17460 28160 17466 28172
rect 18049 28169 18061 28172
rect 18095 28169 18107 28203
rect 22373 28203 22431 28209
rect 18049 28163 18107 28169
rect 18340 28172 22232 28200
rect 11882 28092 11888 28144
rect 11940 28132 11946 28144
rect 12437 28135 12495 28141
rect 12437 28132 12449 28135
rect 11940 28104 12449 28132
rect 11940 28092 11946 28104
rect 12437 28101 12449 28104
rect 12483 28132 12495 28135
rect 13354 28132 13360 28144
rect 12483 28104 13360 28132
rect 12483 28101 12495 28104
rect 12437 28095 12495 28101
rect 13354 28092 13360 28104
rect 13412 28092 13418 28144
rect 14645 28135 14703 28141
rect 14645 28101 14657 28135
rect 14691 28132 14703 28135
rect 18340 28132 18368 28172
rect 14691 28104 18368 28132
rect 18417 28135 18475 28141
rect 14691 28101 14703 28104
rect 14645 28095 14703 28101
rect 18417 28101 18429 28135
rect 18463 28101 18475 28135
rect 18417 28095 18475 28101
rect 18509 28135 18567 28141
rect 18509 28101 18521 28135
rect 18555 28132 18567 28135
rect 18874 28132 18880 28144
rect 18555 28104 18880 28132
rect 18555 28101 18567 28104
rect 18509 28095 18567 28101
rect 12618 28064 12624 28076
rect 10612 28050 12624 28064
rect 10626 28036 12624 28050
rect 9217 28027 9275 28033
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 14090 28024 14096 28076
rect 14148 28064 14154 28076
rect 14274 28064 14280 28076
rect 14148 28036 14280 28064
rect 14148 28024 14154 28036
rect 14274 28024 14280 28036
rect 14332 28064 14338 28076
rect 14737 28067 14795 28073
rect 14737 28064 14749 28067
rect 14332 28036 14749 28064
rect 14332 28024 14338 28036
rect 14737 28033 14749 28036
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28064 17279 28067
rect 18322 28064 18328 28076
rect 17267 28036 18328 28064
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 18322 28024 18328 28036
rect 18380 28024 18386 28076
rect 18432 28008 18460 28095
rect 18874 28092 18880 28104
rect 18932 28092 18938 28144
rect 19797 28135 19855 28141
rect 19797 28101 19809 28135
rect 19843 28132 19855 28135
rect 20530 28132 20536 28144
rect 19843 28104 20536 28132
rect 19843 28101 19855 28104
rect 19797 28095 19855 28101
rect 20530 28092 20536 28104
rect 20588 28092 20594 28144
rect 19337 28067 19395 28073
rect 19337 28064 19349 28067
rect 18708 28036 19349 28064
rect 6270 27956 6276 28008
rect 6328 27996 6334 28008
rect 6549 27999 6607 28005
rect 6549 27996 6561 27999
rect 6328 27968 6561 27996
rect 6328 27956 6334 27968
rect 6549 27965 6561 27968
rect 6595 27965 6607 27999
rect 6549 27959 6607 27965
rect 6825 27999 6883 28005
rect 6825 27965 6837 27999
rect 6871 27996 6883 27999
rect 8294 27996 8300 28008
rect 6871 27968 8300 27996
rect 6871 27965 6883 27968
rect 6825 27959 6883 27965
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27996 9551 27999
rect 10778 27996 10784 28008
rect 9539 27968 10784 27996
rect 9539 27965 9551 27968
rect 9493 27959 9551 27965
rect 10778 27956 10784 27968
rect 10836 27956 10842 28008
rect 12529 27999 12587 28005
rect 12084 27968 12434 27996
rect 10870 27888 10876 27940
rect 10928 27928 10934 27940
rect 11977 27931 12035 27937
rect 11977 27928 11989 27931
rect 10928 27900 11989 27928
rect 10928 27888 10934 27900
rect 11977 27897 11989 27900
rect 12023 27897 12035 27931
rect 11977 27891 12035 27897
rect 7558 27820 7564 27872
rect 7616 27860 7622 27872
rect 12084 27860 12112 27968
rect 12406 27928 12434 27968
rect 12529 27965 12541 27999
rect 12575 27965 12587 27999
rect 12529 27959 12587 27965
rect 14829 27999 14887 28005
rect 14829 27965 14841 27999
rect 14875 27965 14887 27999
rect 14829 27959 14887 27965
rect 12544 27928 12572 27959
rect 14277 27931 14335 27937
rect 14277 27928 14289 27931
rect 12406 27900 12572 27928
rect 12912 27900 14289 27928
rect 7616 27832 12112 27860
rect 7616 27820 7622 27832
rect 12342 27820 12348 27872
rect 12400 27860 12406 27872
rect 12912 27860 12940 27900
rect 14277 27897 14289 27900
rect 14323 27897 14335 27931
rect 14277 27891 14335 27897
rect 14366 27888 14372 27940
rect 14424 27928 14430 27940
rect 14844 27928 14872 27959
rect 16758 27956 16764 28008
rect 16816 27996 16822 28008
rect 17405 27999 17463 28005
rect 17405 27996 17417 27999
rect 16816 27968 17417 27996
rect 16816 27956 16822 27968
rect 17405 27965 17417 27968
rect 17451 27965 17463 27999
rect 17405 27959 17463 27965
rect 18414 27956 18420 28008
rect 18472 27956 18478 28008
rect 18598 27956 18604 28008
rect 18656 27956 18662 28008
rect 14424 27900 14872 27928
rect 14424 27888 14430 27900
rect 15102 27888 15108 27940
rect 15160 27928 15166 27940
rect 18708 27928 18736 28036
rect 19337 28033 19349 28036
rect 19383 28033 19395 28067
rect 19337 28027 19395 28033
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 22204 28064 22232 28172
rect 22373 28169 22385 28203
rect 22419 28200 22431 28203
rect 22554 28200 22560 28212
rect 22419 28172 22560 28200
rect 22419 28169 22431 28172
rect 22373 28163 22431 28169
rect 22554 28160 22560 28172
rect 22612 28160 22618 28212
rect 23658 28092 23664 28144
rect 23716 28132 23722 28144
rect 24673 28135 24731 28141
rect 24673 28132 24685 28135
rect 23716 28104 24685 28132
rect 23716 28092 23722 28104
rect 24673 28101 24685 28104
rect 24719 28101 24731 28135
rect 24673 28095 24731 28101
rect 22830 28064 22836 28076
rect 19484 28036 21588 28064
rect 22204 28036 22836 28064
rect 19484 28024 19490 28036
rect 19242 27956 19248 28008
rect 19300 27996 19306 28008
rect 19889 27999 19947 28005
rect 19889 27996 19901 27999
rect 19300 27968 19901 27996
rect 19300 27956 19306 27968
rect 19889 27965 19901 27968
rect 19935 27965 19947 27999
rect 19889 27959 19947 27965
rect 20070 27956 20076 28008
rect 20128 27956 20134 28008
rect 21560 27996 21588 28036
rect 22830 28024 22836 28036
rect 22888 28024 22894 28076
rect 23474 28024 23480 28076
rect 23532 28024 23538 28076
rect 24026 28024 24032 28076
rect 24084 28064 24090 28076
rect 24121 28067 24179 28073
rect 24121 28064 24133 28067
rect 24084 28036 24133 28064
rect 24084 28024 24090 28036
rect 24121 28033 24133 28036
rect 24167 28033 24179 28067
rect 24121 28027 24179 28033
rect 22465 27999 22523 28005
rect 22465 27996 22477 27999
rect 21560 27968 22477 27996
rect 22465 27965 22477 27968
rect 22511 27965 22523 27999
rect 22465 27959 22523 27965
rect 22649 27999 22707 28005
rect 22649 27965 22661 27999
rect 22695 27996 22707 27999
rect 23750 27996 23756 28008
rect 22695 27968 23756 27996
rect 22695 27965 22707 27968
rect 22649 27959 22707 27965
rect 23750 27956 23756 27968
rect 23808 27956 23814 28008
rect 15160 27900 18736 27928
rect 19153 27931 19211 27937
rect 15160 27888 15166 27900
rect 19153 27897 19165 27931
rect 19199 27928 19211 27931
rect 22094 27928 22100 27940
rect 19199 27900 22100 27928
rect 19199 27897 19211 27900
rect 19153 27891 19211 27897
rect 22094 27888 22100 27900
rect 22152 27888 22158 27940
rect 12400 27832 12940 27860
rect 12400 27820 12406 27832
rect 13354 27820 13360 27872
rect 13412 27820 13418 27872
rect 16574 27820 16580 27872
rect 16632 27860 16638 27872
rect 16853 27863 16911 27869
rect 16853 27860 16865 27863
rect 16632 27832 16865 27860
rect 16632 27820 16638 27832
rect 16853 27829 16865 27832
rect 16899 27829 16911 27863
rect 16853 27823 16911 27829
rect 19429 27863 19487 27869
rect 19429 27829 19441 27863
rect 19475 27860 19487 27863
rect 19886 27860 19892 27872
rect 19475 27832 19892 27860
rect 19475 27829 19487 27832
rect 19429 27823 19487 27829
rect 19886 27820 19892 27832
rect 19944 27820 19950 27872
rect 21910 27820 21916 27872
rect 21968 27860 21974 27872
rect 22005 27863 22063 27869
rect 22005 27860 22017 27863
rect 21968 27832 22017 27860
rect 21968 27820 21974 27832
rect 22005 27829 22017 27832
rect 22051 27829 22063 27863
rect 22005 27823 22063 27829
rect 23290 27820 23296 27872
rect 23348 27820 23354 27872
rect 23934 27820 23940 27872
rect 23992 27820 23998 27872
rect 24210 27820 24216 27872
rect 24268 27860 24274 27872
rect 24765 27863 24823 27869
rect 24765 27860 24777 27863
rect 24268 27832 24777 27860
rect 24268 27820 24274 27832
rect 24765 27829 24777 27832
rect 24811 27829 24823 27863
rect 24765 27823 24823 27829
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 6536 27659 6594 27665
rect 6536 27625 6548 27659
rect 6582 27656 6594 27659
rect 7834 27656 7840 27668
rect 6582 27628 7840 27656
rect 6582 27625 6594 27628
rect 6536 27619 6594 27625
rect 7834 27616 7840 27628
rect 7892 27616 7898 27668
rect 12618 27616 12624 27668
rect 12676 27656 12682 27668
rect 13078 27656 13084 27668
rect 12676 27628 13084 27656
rect 12676 27616 12682 27628
rect 13078 27616 13084 27628
rect 13136 27616 13142 27668
rect 15286 27616 15292 27668
rect 15344 27656 15350 27668
rect 23290 27656 23296 27668
rect 15344 27628 23296 27656
rect 15344 27616 15350 27628
rect 23290 27616 23296 27628
rect 23348 27616 23354 27668
rect 12526 27548 12532 27600
rect 12584 27588 12590 27600
rect 12584 27560 16252 27588
rect 12584 27548 12590 27560
rect 1302 27480 1308 27532
rect 1360 27520 1366 27532
rect 2041 27523 2099 27529
rect 2041 27520 2053 27523
rect 1360 27492 2053 27520
rect 1360 27480 1366 27492
rect 2041 27489 2053 27492
rect 2087 27489 2099 27523
rect 2041 27483 2099 27489
rect 3326 27480 3332 27532
rect 3384 27520 3390 27532
rect 3973 27523 4031 27529
rect 3973 27520 3985 27523
rect 3384 27492 3985 27520
rect 3384 27480 3390 27492
rect 3973 27489 3985 27492
rect 4019 27489 4031 27523
rect 3973 27483 4031 27489
rect 13357 27523 13415 27529
rect 13357 27489 13369 27523
rect 13403 27520 13415 27523
rect 14458 27520 14464 27532
rect 13403 27492 14464 27520
rect 13403 27489 13415 27492
rect 13357 27483 13415 27489
rect 14458 27480 14464 27492
rect 14516 27480 14522 27532
rect 14734 27480 14740 27532
rect 14792 27480 14798 27532
rect 14921 27523 14979 27529
rect 14921 27489 14933 27523
rect 14967 27520 14979 27523
rect 15930 27520 15936 27532
rect 14967 27492 15936 27520
rect 14967 27489 14979 27492
rect 14921 27483 14979 27489
rect 15930 27480 15936 27492
rect 15988 27480 15994 27532
rect 16224 27529 16252 27560
rect 16298 27548 16304 27600
rect 16356 27588 16362 27600
rect 17957 27591 18015 27597
rect 16356 27560 17356 27588
rect 16356 27548 16362 27560
rect 16209 27523 16267 27529
rect 16209 27489 16221 27523
rect 16255 27520 16267 27523
rect 17034 27520 17040 27532
rect 16255 27492 17040 27520
rect 16255 27489 16267 27492
rect 16209 27483 16267 27489
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 17218 27480 17224 27532
rect 17276 27480 17282 27532
rect 17328 27529 17356 27560
rect 17957 27557 17969 27591
rect 18003 27588 18015 27591
rect 19518 27588 19524 27600
rect 18003 27560 19524 27588
rect 18003 27557 18015 27560
rect 17957 27551 18015 27557
rect 19518 27548 19524 27560
rect 19576 27548 19582 27600
rect 23750 27548 23756 27600
rect 23808 27588 23814 27600
rect 24029 27591 24087 27597
rect 24029 27588 24041 27591
rect 23808 27560 24041 27588
rect 23808 27548 23814 27560
rect 24029 27557 24041 27560
rect 24075 27557 24087 27591
rect 24029 27551 24087 27557
rect 17313 27523 17371 27529
rect 17313 27489 17325 27523
rect 17359 27489 17371 27523
rect 17313 27483 17371 27489
rect 18414 27480 18420 27532
rect 18472 27480 18478 27532
rect 18506 27480 18512 27532
rect 18564 27480 18570 27532
rect 22557 27523 22615 27529
rect 22557 27489 22569 27523
rect 22603 27520 22615 27523
rect 23290 27520 23296 27532
rect 22603 27492 23296 27520
rect 22603 27489 22615 27492
rect 22557 27483 22615 27489
rect 23290 27480 23296 27492
rect 23348 27480 23354 27532
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 1946 27452 1952 27464
rect 1811 27424 1952 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 1946 27412 1952 27424
rect 2004 27412 2010 27464
rect 6270 27412 6276 27464
rect 6328 27412 6334 27464
rect 10502 27412 10508 27464
rect 10560 27452 10566 27464
rect 10781 27455 10839 27461
rect 10781 27452 10793 27455
rect 10560 27424 10793 27452
rect 10560 27412 10566 27424
rect 10781 27421 10793 27424
rect 10827 27421 10839 27455
rect 10781 27415 10839 27421
rect 13081 27455 13139 27461
rect 13081 27421 13093 27455
rect 13127 27452 13139 27455
rect 13170 27452 13176 27464
rect 13127 27424 13176 27452
rect 13127 27421 13139 27424
rect 13081 27415 13139 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 16942 27412 16948 27464
rect 17000 27452 17006 27464
rect 17129 27455 17187 27461
rect 17129 27452 17141 27455
rect 17000 27424 17141 27452
rect 17000 27412 17006 27424
rect 17129 27421 17141 27424
rect 17175 27421 17187 27455
rect 17129 27415 17187 27421
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 18012 27424 18337 27452
rect 18012 27412 18018 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 22186 27412 22192 27464
rect 22244 27452 22250 27464
rect 22281 27455 22339 27461
rect 22281 27452 22293 27455
rect 22244 27424 22293 27452
rect 22244 27412 22250 27424
rect 22281 27421 22293 27424
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 23842 27412 23848 27464
rect 23900 27452 23906 27464
rect 24673 27455 24731 27461
rect 24673 27452 24685 27455
rect 23900 27424 24685 27452
rect 23900 27412 23906 27424
rect 24673 27421 24685 27424
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 4157 27387 4215 27393
rect 4157 27384 4169 27387
rect 4080 27356 4169 27384
rect 4080 27328 4108 27356
rect 4157 27353 4169 27356
rect 4203 27353 4215 27387
rect 4157 27347 4215 27353
rect 5813 27387 5871 27393
rect 5813 27353 5825 27387
rect 5859 27384 5871 27387
rect 6086 27384 6092 27396
rect 5859 27356 6092 27384
rect 5859 27353 5871 27356
rect 5813 27347 5871 27353
rect 6086 27344 6092 27356
rect 6144 27344 6150 27396
rect 7282 27344 7288 27396
rect 7340 27344 7346 27396
rect 14645 27387 14703 27393
rect 14645 27384 14657 27387
rect 12728 27356 14657 27384
rect 4062 27276 4068 27328
rect 4120 27276 4126 27328
rect 8021 27319 8079 27325
rect 8021 27285 8033 27319
rect 8067 27316 8079 27319
rect 8386 27316 8392 27328
rect 8067 27288 8392 27316
rect 8067 27285 8079 27288
rect 8021 27279 8079 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 12728 27325 12756 27356
rect 14645 27353 14657 27356
rect 14691 27353 14703 27387
rect 14645 27347 14703 27353
rect 15654 27344 15660 27396
rect 15712 27384 15718 27396
rect 15933 27387 15991 27393
rect 15933 27384 15945 27387
rect 15712 27356 15945 27384
rect 15712 27344 15718 27356
rect 15933 27353 15945 27356
rect 15979 27384 15991 27387
rect 16114 27384 16120 27396
rect 15979 27356 16120 27384
rect 15979 27353 15991 27356
rect 15933 27347 15991 27353
rect 16114 27344 16120 27356
rect 16172 27344 16178 27396
rect 18598 27344 18604 27396
rect 18656 27384 18662 27396
rect 22462 27384 22468 27396
rect 18656 27356 22468 27384
rect 18656 27344 18662 27356
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 24118 27384 24124 27396
rect 23782 27356 24124 27384
rect 24118 27344 24124 27356
rect 24176 27344 24182 27396
rect 24854 27344 24860 27396
rect 24912 27344 24918 27396
rect 12713 27319 12771 27325
rect 12713 27285 12725 27319
rect 12759 27285 12771 27319
rect 12713 27279 12771 27285
rect 13170 27276 13176 27328
rect 13228 27276 13234 27328
rect 13906 27276 13912 27328
rect 13964 27316 13970 27328
rect 14277 27319 14335 27325
rect 14277 27316 14289 27319
rect 13964 27288 14289 27316
rect 13964 27276 13970 27288
rect 14277 27285 14289 27288
rect 14323 27285 14335 27319
rect 14277 27279 14335 27285
rect 15562 27276 15568 27328
rect 15620 27276 15626 27328
rect 16022 27276 16028 27328
rect 16080 27276 16086 27328
rect 16761 27319 16819 27325
rect 16761 27285 16773 27319
rect 16807 27316 16819 27319
rect 17218 27316 17224 27328
rect 16807 27288 17224 27316
rect 16807 27285 16819 27288
rect 16761 27279 16819 27285
rect 17218 27276 17224 27288
rect 17276 27276 17282 27328
rect 17770 27276 17776 27328
rect 17828 27316 17834 27328
rect 23842 27316 23848 27328
rect 17828 27288 23848 27316
rect 17828 27276 17834 27288
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 1762 27072 1768 27124
rect 1820 27112 1826 27124
rect 3510 27121 3516 27124
rect 2041 27115 2099 27121
rect 2041 27112 2053 27115
rect 1820 27084 2053 27112
rect 1820 27072 1826 27084
rect 2041 27081 2053 27084
rect 2087 27081 2099 27115
rect 2041 27075 2099 27081
rect 3467 27115 3516 27121
rect 3467 27081 3479 27115
rect 3513 27081 3516 27115
rect 3467 27075 3516 27081
rect 3510 27072 3516 27075
rect 3568 27072 3574 27124
rect 10410 27072 10416 27124
rect 10468 27072 10474 27124
rect 10778 27072 10784 27124
rect 10836 27112 10842 27124
rect 13449 27115 13507 27121
rect 13449 27112 13461 27115
rect 10836 27084 13461 27112
rect 10836 27072 10842 27084
rect 13449 27081 13461 27084
rect 13495 27112 13507 27115
rect 13998 27112 14004 27124
rect 13495 27084 14004 27112
rect 13495 27081 13507 27084
rect 13449 27075 13507 27081
rect 13998 27072 14004 27084
rect 14056 27072 14062 27124
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 15746 27112 15752 27124
rect 15160 27084 15752 27112
rect 15160 27072 15166 27084
rect 15746 27072 15752 27084
rect 15804 27112 15810 27124
rect 15804 27084 15976 27112
rect 15804 27072 15810 27084
rect 5902 27004 5908 27056
rect 5960 27044 5966 27056
rect 6086 27044 6092 27056
rect 5960 27016 6092 27044
rect 5960 27004 5966 27016
rect 6086 27004 6092 27016
rect 6144 27044 6150 27056
rect 12066 27044 12072 27056
rect 6144 27016 12072 27044
rect 6144 27004 6150 27016
rect 12066 27004 12072 27016
rect 12124 27004 12130 27056
rect 2225 26979 2283 26985
rect 2225 26945 2237 26979
rect 2271 26976 2283 26979
rect 2866 26976 2872 26988
rect 2271 26948 2872 26976
rect 2271 26945 2283 26948
rect 2225 26939 2283 26945
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 3396 26979 3454 26985
rect 3396 26945 3408 26979
rect 3442 26976 3454 26979
rect 3602 26976 3608 26988
rect 3442 26948 3608 26976
rect 3442 26945 3454 26948
rect 3396 26939 3454 26945
rect 3602 26936 3608 26948
rect 3660 26936 3666 26988
rect 7929 26979 7987 26985
rect 7929 26945 7941 26979
rect 7975 26976 7987 26979
rect 9306 26976 9312 26988
rect 7975 26948 9312 26976
rect 7975 26945 7987 26948
rect 7929 26939 7987 26945
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 10321 26979 10379 26985
rect 10321 26976 10333 26979
rect 9456 26948 10333 26976
rect 9456 26936 9462 26948
rect 10321 26945 10333 26948
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 11238 26936 11244 26988
rect 11296 26976 11302 26988
rect 11422 26976 11428 26988
rect 11296 26948 11428 26976
rect 11296 26936 11302 26948
rect 11422 26936 11428 26948
rect 11480 26976 11486 26988
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11480 26948 11713 26976
rect 11480 26936 11486 26948
rect 11701 26945 11713 26948
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 13078 26936 13084 26988
rect 13136 26976 13142 26988
rect 13998 26976 14004 26988
rect 13136 26948 14004 26976
rect 13136 26936 13142 26948
rect 13998 26936 14004 26948
rect 14056 26936 14062 26988
rect 14090 26936 14096 26988
rect 14148 26976 14154 26988
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14148 26948 15025 26976
rect 14148 26936 14154 26948
rect 15013 26945 15025 26948
rect 15059 26976 15071 26979
rect 15948 26976 15976 27084
rect 17494 27072 17500 27124
rect 17552 27112 17558 27124
rect 17862 27112 17868 27124
rect 17552 27084 17868 27112
rect 17552 27072 17558 27084
rect 17862 27072 17868 27084
rect 17920 27072 17926 27124
rect 20346 27112 20352 27124
rect 19352 27084 20352 27112
rect 16022 27004 16028 27056
rect 16080 27044 16086 27056
rect 18782 27044 18788 27056
rect 16080 27016 18788 27044
rect 16080 27004 16086 27016
rect 18782 27004 18788 27016
rect 18840 27004 18846 27056
rect 19352 26985 19380 27084
rect 20346 27072 20352 27084
rect 20404 27112 20410 27124
rect 22186 27112 22192 27124
rect 20404 27084 22192 27112
rect 20404 27072 20410 27084
rect 22186 27072 22192 27084
rect 22244 27072 22250 27124
rect 22462 27072 22468 27124
rect 22520 27112 22526 27124
rect 23937 27115 23995 27121
rect 23937 27112 23949 27115
rect 22520 27084 23949 27112
rect 22520 27072 22526 27084
rect 23937 27081 23949 27084
rect 23983 27081 23995 27115
rect 23937 27075 23995 27081
rect 19610 27004 19616 27056
rect 19668 27004 19674 27056
rect 21266 27044 21272 27056
rect 20838 27016 21272 27044
rect 21266 27004 21272 27016
rect 21324 27004 21330 27056
rect 24118 27044 24124 27056
rect 23690 27016 24124 27044
rect 24118 27004 24124 27016
rect 24176 27004 24182 27056
rect 24670 27004 24676 27056
rect 24728 27004 24734 27056
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 15059 26948 15792 26976
rect 15948 26948 17785 26976
rect 15059 26945 15071 26948
rect 15013 26939 15071 26945
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 8021 26911 8079 26917
rect 8021 26908 8033 26911
rect 7432 26880 8033 26908
rect 7432 26868 7438 26880
rect 8021 26877 8033 26880
rect 8067 26877 8079 26911
rect 8021 26871 8079 26877
rect 8113 26911 8171 26917
rect 8113 26877 8125 26911
rect 8159 26877 8171 26911
rect 8113 26871 8171 26877
rect 7742 26840 7748 26852
rect 6886 26812 7748 26840
rect 4890 26732 4896 26784
rect 4948 26772 4954 26784
rect 6886 26772 6914 26812
rect 7742 26800 7748 26812
rect 7800 26800 7806 26852
rect 7834 26800 7840 26852
rect 7892 26840 7898 26852
rect 8128 26840 8156 26871
rect 8294 26868 8300 26920
rect 8352 26908 8358 26920
rect 10505 26911 10563 26917
rect 10505 26908 10517 26911
rect 8352 26880 10517 26908
rect 8352 26868 8358 26880
rect 10505 26877 10517 26880
rect 10551 26877 10563 26911
rect 10505 26871 10563 26877
rect 11977 26911 12035 26917
rect 11977 26877 11989 26911
rect 12023 26908 12035 26911
rect 13446 26908 13452 26920
rect 12023 26880 13452 26908
rect 12023 26877 12035 26880
rect 11977 26871 12035 26877
rect 13446 26868 13452 26880
rect 13504 26868 13510 26920
rect 15102 26868 15108 26920
rect 15160 26868 15166 26920
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26877 15255 26911
rect 15764 26908 15792 26948
rect 17773 26945 17785 26948
rect 17819 26945 17831 26979
rect 19337 26979 19395 26985
rect 17773 26939 17831 26945
rect 17972 26948 19288 26976
rect 17972 26908 18000 26948
rect 15764 26880 18000 26908
rect 18049 26911 18107 26917
rect 15197 26871 15255 26877
rect 18049 26877 18061 26911
rect 18095 26908 18107 26911
rect 18690 26908 18696 26920
rect 18095 26880 18696 26908
rect 18095 26877 18107 26880
rect 18049 26871 18107 26877
rect 7892 26812 8156 26840
rect 7892 26800 7898 26812
rect 12986 26800 12992 26852
rect 13044 26840 13050 26852
rect 15212 26840 15240 26871
rect 13044 26812 15240 26840
rect 13044 26800 13050 26812
rect 17126 26800 17132 26852
rect 17184 26840 17190 26852
rect 18064 26840 18092 26871
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 19260 26908 19288 26948
rect 19337 26945 19349 26979
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19702 26908 19708 26920
rect 19260 26880 19708 26908
rect 19702 26868 19708 26880
rect 19760 26868 19766 26920
rect 20070 26868 20076 26920
rect 20128 26908 20134 26920
rect 20622 26908 20628 26920
rect 20128 26880 20628 26908
rect 20128 26868 20134 26880
rect 20622 26868 20628 26880
rect 20680 26908 20686 26920
rect 21085 26911 21143 26917
rect 21085 26908 21097 26911
rect 20680 26880 21097 26908
rect 20680 26868 20686 26880
rect 21085 26877 21097 26880
rect 21131 26877 21143 26911
rect 21085 26871 21143 26877
rect 22186 26868 22192 26920
rect 22244 26868 22250 26920
rect 22462 26868 22468 26920
rect 22520 26868 22526 26920
rect 17184 26812 18092 26840
rect 17184 26800 17190 26812
rect 4948 26744 6914 26772
rect 4948 26732 4954 26744
rect 7006 26732 7012 26784
rect 7064 26772 7070 26784
rect 7282 26772 7288 26784
rect 7064 26744 7288 26772
rect 7064 26732 7070 26744
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 7561 26775 7619 26781
rect 7561 26741 7573 26775
rect 7607 26772 7619 26775
rect 8570 26772 8576 26784
rect 7607 26744 8576 26772
rect 7607 26741 7619 26744
rect 7561 26735 7619 26741
rect 8570 26732 8576 26744
rect 8628 26732 8634 26784
rect 8938 26732 8944 26784
rect 8996 26732 9002 26784
rect 9953 26775 10011 26781
rect 9953 26741 9965 26775
rect 9999 26772 10011 26775
rect 11974 26772 11980 26784
rect 9999 26744 11980 26772
rect 9999 26741 10011 26744
rect 9953 26735 10011 26741
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 14642 26732 14648 26784
rect 14700 26732 14706 26784
rect 17402 26732 17408 26784
rect 17460 26732 17466 26784
rect 20254 26732 20260 26784
rect 20312 26772 20318 26784
rect 23198 26772 23204 26784
rect 20312 26744 23204 26772
rect 20312 26732 20318 26744
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 24765 26775 24823 26781
rect 24765 26772 24777 26775
rect 23624 26744 24777 26772
rect 23624 26732 23630 26744
rect 24765 26741 24777 26744
rect 24811 26741 24823 26775
rect 24765 26735 24823 26741
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 7098 26528 7104 26580
rect 7156 26568 7162 26580
rect 7558 26568 7564 26580
rect 7156 26540 7564 26568
rect 7156 26528 7162 26540
rect 7558 26528 7564 26540
rect 7616 26568 7622 26580
rect 8021 26571 8079 26577
rect 8021 26568 8033 26571
rect 7616 26540 8033 26568
rect 7616 26528 7622 26540
rect 8021 26537 8033 26540
rect 8067 26537 8079 26571
rect 8021 26531 8079 26537
rect 9306 26528 9312 26580
rect 9364 26528 9370 26580
rect 11054 26528 11060 26580
rect 11112 26568 11118 26580
rect 11112 26540 11744 26568
rect 11112 26528 11118 26540
rect 7742 26460 7748 26512
rect 7800 26500 7806 26512
rect 10042 26500 10048 26512
rect 7800 26472 10048 26500
rect 7800 26460 7806 26472
rect 10042 26460 10048 26472
rect 10100 26460 10106 26512
rect 10137 26503 10195 26509
rect 10137 26469 10149 26503
rect 10183 26500 10195 26503
rect 10183 26472 11652 26500
rect 10183 26469 10195 26472
rect 10137 26463 10195 26469
rect 1578 26392 1584 26444
rect 1636 26432 1642 26444
rect 3973 26435 4031 26441
rect 3973 26432 3985 26435
rect 1636 26404 3985 26432
rect 1636 26392 1642 26404
rect 3973 26401 3985 26404
rect 4019 26401 4031 26435
rect 3973 26395 4031 26401
rect 4890 26392 4896 26444
rect 4948 26392 4954 26444
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 6595 26404 7788 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 7760 26364 7788 26404
rect 10778 26392 10784 26444
rect 10836 26392 10842 26444
rect 8386 26364 8392 26376
rect 7760 26336 8392 26364
rect 8386 26324 8392 26336
rect 8444 26324 8450 26376
rect 10502 26324 10508 26376
rect 10560 26324 10566 26376
rect 11624 26364 11652 26472
rect 11716 26432 11744 26540
rect 13170 26528 13176 26580
rect 13228 26568 13234 26580
rect 13998 26568 14004 26580
rect 13228 26540 14004 26568
rect 13228 26528 13234 26540
rect 13998 26528 14004 26540
rect 14056 26568 14062 26580
rect 15378 26568 15384 26580
rect 14056 26540 15384 26568
rect 14056 26528 14062 26540
rect 15378 26528 15384 26540
rect 15436 26568 15442 26580
rect 16022 26568 16028 26580
rect 15436 26540 16028 26568
rect 15436 26528 15442 26540
rect 16022 26528 16028 26540
rect 16080 26528 16086 26580
rect 16206 26528 16212 26580
rect 16264 26568 16270 26580
rect 16758 26568 16764 26580
rect 16264 26540 16764 26568
rect 16264 26528 16270 26540
rect 16758 26528 16764 26540
rect 16816 26528 16822 26580
rect 19797 26571 19855 26577
rect 19797 26537 19809 26571
rect 19843 26568 19855 26571
rect 22370 26568 22376 26580
rect 19843 26540 22376 26568
rect 19843 26537 19855 26540
rect 19797 26531 19855 26537
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 23201 26571 23259 26577
rect 23201 26537 23213 26571
rect 23247 26568 23259 26571
rect 23290 26568 23296 26580
rect 23247 26540 23296 26568
rect 23247 26537 23259 26540
rect 23201 26531 23259 26537
rect 23290 26528 23296 26540
rect 23348 26528 23354 26580
rect 23842 26528 23848 26580
rect 23900 26528 23906 26580
rect 12713 26503 12771 26509
rect 12713 26469 12725 26503
rect 12759 26500 12771 26503
rect 13722 26500 13728 26512
rect 12759 26472 13728 26500
rect 12759 26469 12771 26472
rect 12713 26463 12771 26469
rect 13722 26460 13728 26472
rect 13780 26460 13786 26512
rect 13265 26435 13323 26441
rect 13265 26432 13277 26435
rect 11716 26404 13277 26432
rect 13265 26401 13277 26404
rect 13311 26401 13323 26435
rect 13265 26395 13323 26401
rect 14182 26392 14188 26444
rect 14240 26432 14246 26444
rect 17770 26432 17776 26444
rect 14240 26404 17776 26432
rect 14240 26392 14246 26404
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 20254 26392 20260 26444
rect 20312 26432 20318 26444
rect 20349 26435 20407 26441
rect 20349 26432 20361 26435
rect 20312 26404 20361 26432
rect 20312 26392 20318 26404
rect 20349 26401 20361 26404
rect 20395 26401 20407 26435
rect 20349 26395 20407 26401
rect 21453 26435 21511 26441
rect 21453 26401 21465 26435
rect 21499 26432 21511 26435
rect 22186 26432 22192 26444
rect 21499 26404 22192 26432
rect 21499 26401 21511 26404
rect 21453 26395 21511 26401
rect 22186 26392 22192 26404
rect 22244 26432 22250 26444
rect 22738 26432 22744 26444
rect 22244 26404 22744 26432
rect 22244 26392 22250 26404
rect 22738 26392 22744 26404
rect 22796 26392 22802 26444
rect 13081 26367 13139 26373
rect 13081 26364 13093 26367
rect 11624 26336 13093 26364
rect 13081 26333 13093 26336
rect 13127 26333 13139 26367
rect 13081 26327 13139 26333
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26364 13231 26367
rect 13538 26364 13544 26376
rect 13219 26336 13544 26364
rect 13219 26333 13231 26336
rect 13173 26327 13231 26333
rect 13538 26324 13544 26336
rect 13596 26324 13602 26376
rect 14458 26324 14464 26376
rect 14516 26324 14522 26376
rect 24029 26367 24087 26373
rect 24029 26333 24041 26367
rect 24075 26364 24087 26367
rect 24946 26364 24952 26376
rect 24075 26336 24952 26364
rect 24075 26333 24087 26336
rect 24029 26327 24087 26333
rect 24946 26324 24952 26336
rect 25004 26324 25010 26376
rect 3878 26256 3884 26308
rect 3936 26296 3942 26308
rect 4157 26299 4215 26305
rect 4157 26296 4169 26299
rect 3936 26268 4169 26296
rect 3936 26256 3942 26268
rect 4157 26265 4169 26268
rect 4203 26265 4215 26299
rect 6288 26296 6316 26324
rect 6454 26296 6460 26308
rect 6288 26268 6460 26296
rect 4157 26259 4215 26265
rect 6454 26256 6460 26268
rect 6512 26256 6518 26308
rect 7282 26256 7288 26308
rect 7340 26256 7346 26308
rect 10594 26256 10600 26308
rect 10652 26256 10658 26308
rect 14737 26299 14795 26305
rect 14737 26265 14749 26299
rect 14783 26296 14795 26299
rect 16022 26296 16028 26308
rect 14783 26268 15148 26296
rect 15962 26268 16028 26296
rect 14783 26265 14795 26268
rect 14737 26259 14795 26265
rect 15120 26228 15148 26268
rect 16022 26256 16028 26268
rect 16080 26256 16086 26308
rect 16850 26296 16856 26308
rect 16408 26268 16856 26296
rect 16408 26240 16436 26268
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 19978 26256 19984 26308
rect 20036 26296 20042 26308
rect 20257 26299 20315 26305
rect 20257 26296 20269 26299
rect 20036 26268 20269 26296
rect 20036 26256 20042 26268
rect 20257 26265 20269 26268
rect 20303 26265 20315 26299
rect 20257 26259 20315 26265
rect 21634 26256 21640 26308
rect 21692 26296 21698 26308
rect 21729 26299 21787 26305
rect 21729 26296 21741 26299
rect 21692 26268 21741 26296
rect 21692 26256 21698 26268
rect 21729 26265 21741 26268
rect 21775 26265 21787 26299
rect 24118 26296 24124 26308
rect 22954 26268 24124 26296
rect 21729 26259 21787 26265
rect 16390 26228 16396 26240
rect 15120 26200 16396 26228
rect 16390 26188 16396 26200
rect 16448 26188 16454 26240
rect 16758 26188 16764 26240
rect 16816 26228 16822 26240
rect 17310 26228 17316 26240
rect 16816 26200 17316 26228
rect 16816 26188 16822 26200
rect 17310 26188 17316 26200
rect 17368 26228 17374 26240
rect 20165 26231 20223 26237
rect 20165 26228 20177 26231
rect 17368 26200 20177 26228
rect 17368 26188 17374 26200
rect 20165 26197 20177 26200
rect 20211 26197 20223 26231
rect 20165 26191 20223 26197
rect 21266 26188 21272 26240
rect 21324 26228 21330 26240
rect 23032 26228 23060 26268
rect 24118 26256 24124 26268
rect 24176 26256 24182 26308
rect 24302 26256 24308 26308
rect 24360 26296 24366 26308
rect 24673 26299 24731 26305
rect 24673 26296 24685 26299
rect 24360 26268 24685 26296
rect 24360 26256 24366 26268
rect 24673 26265 24685 26268
rect 24719 26265 24731 26299
rect 24673 26259 24731 26265
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 25038 26296 25044 26308
rect 24903 26268 25044 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 21324 26200 23060 26228
rect 21324 26188 21330 26200
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 3835 26027 3893 26033
rect 3835 25993 3847 26027
rect 3881 26024 3893 26027
rect 3970 26024 3976 26036
rect 3881 25996 3976 26024
rect 3881 25993 3893 25996
rect 3835 25987 3893 25993
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 26024 7895 26027
rect 8938 26024 8944 26036
rect 7883 25996 8944 26024
rect 7883 25993 7895 25996
rect 7837 25987 7895 25993
rect 8938 25984 8944 25996
rect 8996 25984 9002 26036
rect 10226 25984 10232 26036
rect 10284 26024 10290 26036
rect 10413 26027 10471 26033
rect 10413 26024 10425 26027
rect 10284 25996 10425 26024
rect 10284 25984 10290 25996
rect 10413 25993 10425 25996
rect 10459 25993 10471 26027
rect 10413 25987 10471 25993
rect 15286 25984 15292 26036
rect 15344 26024 15350 26036
rect 16025 26027 16083 26033
rect 16025 26024 16037 26027
rect 15344 25996 16037 26024
rect 15344 25984 15350 25996
rect 16025 25993 16037 25996
rect 16071 25993 16083 26027
rect 16025 25987 16083 25993
rect 17405 26027 17463 26033
rect 17405 25993 17417 26027
rect 17451 26024 17463 26027
rect 19426 26024 19432 26036
rect 17451 25996 19432 26024
rect 17451 25993 17463 25996
rect 17405 25987 17463 25993
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 19518 25984 19524 26036
rect 19576 25984 19582 26036
rect 21082 25984 21088 26036
rect 21140 26024 21146 26036
rect 21269 26027 21327 26033
rect 21269 26024 21281 26027
rect 21140 25996 21281 26024
rect 21140 25984 21146 25996
rect 21269 25993 21281 25996
rect 21315 25993 21327 26027
rect 21269 25987 21327 25993
rect 22002 25984 22008 26036
rect 22060 26024 22066 26036
rect 22060 25984 22094 26024
rect 22278 25984 22284 26036
rect 22336 26024 22342 26036
rect 22373 26027 22431 26033
rect 22373 26024 22385 26027
rect 22336 25996 22385 26024
rect 22336 25984 22342 25996
rect 22373 25993 22385 25996
rect 22419 26024 22431 26027
rect 23201 26027 23259 26033
rect 23201 26024 23213 26027
rect 22419 25996 23213 26024
rect 22419 25993 22431 25996
rect 22373 25987 22431 25993
rect 23201 25993 23213 25996
rect 23247 25993 23259 26027
rect 23201 25987 23259 25993
rect 8570 25916 8576 25968
rect 8628 25956 8634 25968
rect 10321 25959 10379 25965
rect 10321 25956 10333 25959
rect 8628 25928 10333 25956
rect 8628 25916 8634 25928
rect 10321 25925 10333 25928
rect 10367 25925 10379 25959
rect 10321 25919 10379 25925
rect 15102 25916 15108 25968
rect 15160 25956 15166 25968
rect 15933 25959 15991 25965
rect 15933 25956 15945 25959
rect 15160 25928 15945 25956
rect 15160 25916 15166 25928
rect 15933 25925 15945 25928
rect 15979 25956 15991 25959
rect 16758 25956 16764 25968
rect 15979 25928 16764 25956
rect 15979 25925 15991 25928
rect 15933 25919 15991 25925
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25956 17831 25959
rect 17862 25956 17868 25968
rect 17819 25928 17868 25956
rect 17819 25925 17831 25928
rect 17773 25919 17831 25925
rect 17862 25916 17868 25928
rect 17920 25916 17926 25968
rect 22066 25956 22094 25984
rect 24213 25959 24271 25965
rect 24213 25956 24225 25959
rect 22066 25928 24225 25956
rect 24213 25925 24225 25928
rect 24259 25925 24271 25959
rect 24213 25919 24271 25925
rect 24949 25959 25007 25965
rect 24949 25925 24961 25959
rect 24995 25956 25007 25959
rect 25222 25956 25228 25968
rect 24995 25928 25228 25956
rect 24995 25925 25007 25928
rect 24949 25919 25007 25925
rect 25222 25916 25228 25928
rect 25280 25916 25286 25968
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 3326 25888 3332 25900
rect 2639 25860 3332 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 3326 25848 3332 25860
rect 3384 25848 3390 25900
rect 3418 25848 3424 25900
rect 3476 25888 3482 25900
rect 3732 25891 3790 25897
rect 3732 25888 3744 25891
rect 3476 25860 3744 25888
rect 3476 25848 3482 25860
rect 3732 25857 3744 25860
rect 3778 25857 3790 25891
rect 3732 25851 3790 25857
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 6972 25860 8064 25888
rect 6972 25848 6978 25860
rect 2777 25823 2835 25829
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 3602 25820 3608 25832
rect 2823 25792 3608 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 7190 25820 7196 25832
rect 6886 25792 7196 25820
rect 2866 25712 2872 25764
rect 2924 25752 2930 25764
rect 2961 25755 3019 25761
rect 2961 25752 2973 25755
rect 2924 25724 2973 25752
rect 2924 25712 2930 25724
rect 2961 25721 2973 25724
rect 3007 25721 3019 25755
rect 2961 25715 3019 25721
rect 3786 25712 3792 25764
rect 3844 25752 3850 25764
rect 6886 25752 6914 25792
rect 7190 25780 7196 25792
rect 7248 25820 7254 25832
rect 8036 25829 8064 25860
rect 13170 25848 13176 25900
rect 13228 25848 13234 25900
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25888 19487 25891
rect 20438 25888 20444 25900
rect 19475 25860 20444 25888
rect 19475 25857 19487 25860
rect 19429 25851 19487 25857
rect 20438 25848 20444 25860
rect 20496 25848 20502 25900
rect 21453 25891 21511 25897
rect 21453 25857 21465 25891
rect 21499 25888 21511 25891
rect 22278 25888 22284 25900
rect 21499 25860 22284 25888
rect 21499 25857 21511 25860
rect 21453 25851 21511 25857
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 23477 25891 23535 25897
rect 23477 25888 23489 25891
rect 22388 25860 23489 25888
rect 7929 25823 7987 25829
rect 7929 25820 7941 25823
rect 7248 25792 7941 25820
rect 7248 25780 7254 25792
rect 7929 25789 7941 25792
rect 7975 25789 7987 25823
rect 7929 25783 7987 25789
rect 8021 25823 8079 25829
rect 8021 25789 8033 25823
rect 8067 25789 8079 25823
rect 8021 25783 8079 25789
rect 8386 25780 8392 25832
rect 8444 25820 8450 25832
rect 10505 25823 10563 25829
rect 10505 25820 10517 25823
rect 8444 25792 10517 25820
rect 8444 25780 8450 25792
rect 10505 25789 10517 25792
rect 10551 25789 10563 25823
rect 10505 25783 10563 25789
rect 11422 25780 11428 25832
rect 11480 25820 11486 25832
rect 11790 25820 11796 25832
rect 11480 25792 11796 25820
rect 11480 25780 11486 25792
rect 11790 25780 11796 25792
rect 11848 25780 11854 25832
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25820 12127 25823
rect 12802 25820 12808 25832
rect 12115 25792 12808 25820
rect 12115 25789 12127 25792
rect 12069 25783 12127 25789
rect 12802 25780 12808 25792
rect 12860 25780 12866 25832
rect 16209 25823 16267 25829
rect 16209 25789 16221 25823
rect 16255 25820 16267 25823
rect 16390 25820 16396 25832
rect 16255 25792 16396 25820
rect 16255 25789 16267 25792
rect 16209 25783 16267 25789
rect 16390 25780 16396 25792
rect 16448 25780 16454 25832
rect 17770 25780 17776 25832
rect 17828 25820 17834 25832
rect 17865 25823 17923 25829
rect 17865 25820 17877 25823
rect 17828 25792 17877 25820
rect 17828 25780 17834 25792
rect 17865 25789 17877 25792
rect 17911 25789 17923 25823
rect 17865 25783 17923 25789
rect 18049 25823 18107 25829
rect 18049 25789 18061 25823
rect 18095 25820 18107 25823
rect 19610 25820 19616 25832
rect 18095 25792 19616 25820
rect 18095 25789 18107 25792
rect 18049 25783 18107 25789
rect 19610 25780 19616 25792
rect 19668 25780 19674 25832
rect 19702 25780 19708 25832
rect 19760 25780 19766 25832
rect 21726 25780 21732 25832
rect 21784 25820 21790 25832
rect 22388 25820 22416 25860
rect 23477 25857 23489 25860
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 21784 25792 22416 25820
rect 22465 25823 22523 25829
rect 21784 25780 21790 25792
rect 22465 25789 22477 25823
rect 22511 25820 22523 25823
rect 22649 25823 22707 25829
rect 22511 25792 22600 25820
rect 22511 25789 22523 25792
rect 22465 25783 22523 25789
rect 3844 25724 6914 25752
rect 7469 25755 7527 25761
rect 3844 25712 3850 25724
rect 7469 25721 7481 25755
rect 7515 25752 7527 25755
rect 9398 25752 9404 25764
rect 7515 25724 9404 25752
rect 7515 25721 7527 25724
rect 7469 25715 7527 25721
rect 9398 25712 9404 25724
rect 9456 25712 9462 25764
rect 10594 25752 10600 25764
rect 9508 25724 10600 25752
rect 7190 25644 7196 25696
rect 7248 25684 7254 25696
rect 9508 25684 9536 25724
rect 10594 25712 10600 25724
rect 10652 25712 10658 25764
rect 13464 25724 13676 25752
rect 7248 25656 9536 25684
rect 9953 25687 10011 25693
rect 7248 25644 7254 25656
rect 9953 25653 9965 25687
rect 9999 25684 10011 25687
rect 13464 25684 13492 25724
rect 9999 25656 13492 25684
rect 9999 25653 10011 25656
rect 9953 25647 10011 25653
rect 13538 25644 13544 25696
rect 13596 25644 13602 25696
rect 13648 25684 13676 25724
rect 14550 25712 14556 25764
rect 14608 25752 14614 25764
rect 21450 25752 21456 25764
rect 14608 25724 21456 25752
rect 14608 25712 14614 25724
rect 21450 25712 21456 25724
rect 21508 25712 21514 25764
rect 14918 25684 14924 25696
rect 13648 25656 14924 25684
rect 14918 25644 14924 25656
rect 14976 25644 14982 25696
rect 15565 25687 15623 25693
rect 15565 25653 15577 25687
rect 15611 25684 15623 25687
rect 15746 25684 15752 25696
rect 15611 25656 15752 25684
rect 15611 25653 15623 25656
rect 15565 25647 15623 25653
rect 15746 25644 15752 25656
rect 15804 25644 15810 25696
rect 18690 25644 18696 25696
rect 18748 25684 18754 25696
rect 19061 25687 19119 25693
rect 19061 25684 19073 25687
rect 18748 25656 19073 25684
rect 18748 25644 18754 25656
rect 19061 25653 19073 25656
rect 19107 25653 19119 25687
rect 19061 25647 19119 25653
rect 19518 25644 19524 25696
rect 19576 25684 19582 25696
rect 20441 25687 20499 25693
rect 20441 25684 20453 25687
rect 19576 25656 20453 25684
rect 19576 25644 19582 25656
rect 20441 25653 20453 25656
rect 20487 25653 20499 25687
rect 20441 25647 20499 25653
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21784 25656 22017 25684
rect 21784 25644 21790 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 22572 25684 22600 25792
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 23290 25820 23296 25832
rect 22695 25792 23296 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 23290 25780 23296 25792
rect 23348 25780 23354 25832
rect 23474 25712 23480 25764
rect 23532 25752 23538 25764
rect 23661 25755 23719 25761
rect 23661 25752 23673 25755
rect 23532 25724 23673 25752
rect 23532 25712 23538 25724
rect 23661 25721 23673 25724
rect 23707 25721 23719 25755
rect 23661 25715 23719 25721
rect 25133 25755 25191 25761
rect 25133 25721 25145 25755
rect 25179 25752 25191 25755
rect 25222 25752 25228 25764
rect 25179 25724 25228 25752
rect 25179 25721 25191 25724
rect 25133 25715 25191 25721
rect 25222 25712 25228 25724
rect 25280 25712 25286 25764
rect 22152 25656 22600 25684
rect 22152 25644 22158 25656
rect 22738 25644 22744 25696
rect 22796 25684 22802 25696
rect 24305 25687 24363 25693
rect 24305 25684 24317 25687
rect 22796 25656 24317 25684
rect 22796 25644 22802 25656
rect 24305 25653 24317 25656
rect 24351 25653 24363 25687
rect 24305 25647 24363 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 4249 25483 4307 25489
rect 4249 25449 4261 25483
rect 4295 25480 4307 25483
rect 4614 25480 4620 25492
rect 4295 25452 4620 25480
rect 4295 25449 4307 25452
rect 4249 25443 4307 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 5810 25440 5816 25492
rect 5868 25480 5874 25492
rect 6270 25480 6276 25492
rect 5868 25452 6276 25480
rect 5868 25440 5874 25452
rect 6270 25440 6276 25452
rect 6328 25480 6334 25492
rect 15102 25480 15108 25492
rect 6328 25452 15108 25480
rect 6328 25440 6334 25452
rect 15102 25440 15108 25452
rect 15160 25440 15166 25492
rect 18601 25483 18659 25489
rect 18601 25449 18613 25483
rect 18647 25480 18659 25483
rect 19610 25480 19616 25492
rect 18647 25452 19616 25480
rect 18647 25449 18659 25452
rect 18601 25443 18659 25449
rect 19610 25440 19616 25452
rect 19668 25440 19674 25492
rect 19794 25440 19800 25492
rect 19852 25480 19858 25492
rect 19852 25452 22094 25480
rect 19852 25440 19858 25452
rect 12161 25415 12219 25421
rect 12161 25381 12173 25415
rect 12207 25412 12219 25415
rect 14550 25412 14556 25424
rect 12207 25384 14556 25412
rect 12207 25381 12219 25384
rect 12161 25375 12219 25381
rect 14550 25372 14556 25384
rect 14608 25372 14614 25424
rect 1302 25304 1308 25356
rect 1360 25344 1366 25356
rect 2041 25347 2099 25353
rect 2041 25344 2053 25347
rect 1360 25316 2053 25344
rect 1360 25304 1366 25316
rect 2041 25313 2053 25316
rect 2087 25313 2099 25347
rect 2041 25307 2099 25313
rect 6454 25304 6460 25356
rect 6512 25304 6518 25356
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25344 6791 25347
rect 7098 25344 7104 25356
rect 6779 25316 7104 25344
rect 6779 25313 6791 25316
rect 6733 25307 6791 25313
rect 7098 25304 7104 25316
rect 7156 25344 7162 25356
rect 7466 25344 7472 25356
rect 7156 25316 7472 25344
rect 7156 25304 7162 25316
rect 7466 25304 7472 25316
rect 7524 25304 7530 25356
rect 12802 25304 12808 25356
rect 12860 25304 12866 25356
rect 15562 25304 15568 25356
rect 15620 25304 15626 25356
rect 15654 25304 15660 25356
rect 15712 25304 15718 25356
rect 18322 25304 18328 25356
rect 18380 25344 18386 25356
rect 18380 25316 19656 25344
rect 18380 25304 18386 25316
rect 1762 25236 1768 25288
rect 1820 25236 1826 25288
rect 3694 25236 3700 25288
rect 3752 25276 3758 25288
rect 3970 25276 3976 25288
rect 3752 25248 3976 25276
rect 3752 25236 3758 25248
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 7834 25236 7840 25288
rect 7892 25236 7898 25288
rect 9030 25236 9036 25288
rect 9088 25276 9094 25288
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 9088 25248 9321 25276
rect 9088 25236 9094 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 11330 25276 11336 25288
rect 10551 25248 11336 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25276 12587 25279
rect 13541 25279 13599 25285
rect 13541 25276 13553 25279
rect 12575 25248 13553 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 13541 25245 13553 25248
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 16850 25276 16856 25288
rect 14516 25248 16856 25276
rect 14516 25236 14522 25248
rect 16850 25236 16856 25248
rect 16908 25236 16914 25288
rect 19628 25285 19656 25316
rect 20346 25304 20352 25356
rect 20404 25304 20410 25356
rect 20622 25304 20628 25356
rect 20680 25304 20686 25356
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25245 19671 25279
rect 22066 25276 22094 25452
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 23017 25347 23075 25353
rect 23017 25344 23029 25347
rect 22704 25316 23029 25344
rect 22704 25304 22710 25316
rect 23017 25313 23029 25316
rect 23063 25313 23075 25347
rect 23017 25307 23075 25313
rect 23201 25347 23259 25353
rect 23201 25313 23213 25347
rect 23247 25344 23259 25347
rect 23382 25344 23388 25356
rect 23247 25316 23388 25344
rect 23247 25313 23259 25316
rect 23201 25307 23259 25313
rect 23382 25304 23388 25316
rect 23440 25304 23446 25356
rect 23845 25279 23903 25285
rect 23845 25276 23857 25279
rect 22066 25248 23857 25276
rect 19613 25239 19671 25245
rect 23845 25245 23857 25248
rect 23891 25245 23903 25279
rect 23845 25239 23903 25245
rect 23934 25236 23940 25288
rect 23992 25276 23998 25288
rect 24765 25279 24823 25285
rect 24765 25276 24777 25279
rect 23992 25248 24777 25276
rect 23992 25236 23998 25248
rect 24765 25245 24777 25248
rect 24811 25245 24823 25279
rect 24765 25239 24823 25245
rect 12621 25211 12679 25217
rect 12621 25208 12633 25211
rect 12406 25180 12633 25208
rect 3602 25100 3608 25152
rect 3660 25140 3666 25152
rect 4433 25143 4491 25149
rect 4433 25140 4445 25143
rect 3660 25112 4445 25140
rect 3660 25100 3666 25112
rect 4433 25109 4445 25112
rect 4479 25109 4491 25143
rect 4433 25103 4491 25109
rect 8202 25100 8208 25152
rect 8260 25100 8266 25152
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 10597 25143 10655 25149
rect 10597 25140 10609 25143
rect 9824 25112 10609 25140
rect 9824 25100 9830 25112
rect 10597 25109 10609 25112
rect 10643 25109 10655 25143
rect 10597 25103 10655 25109
rect 11698 25100 11704 25152
rect 11756 25140 11762 25152
rect 12406 25140 12434 25180
rect 12621 25177 12633 25180
rect 12667 25177 12679 25211
rect 12621 25171 12679 25177
rect 16298 25168 16304 25220
rect 16356 25208 16362 25220
rect 17129 25211 17187 25217
rect 17129 25208 17141 25211
rect 16356 25180 17141 25208
rect 16356 25168 16362 25180
rect 17129 25177 17141 25180
rect 17175 25177 17187 25211
rect 19058 25208 19064 25220
rect 18354 25180 19064 25208
rect 17129 25171 17187 25177
rect 19058 25168 19064 25180
rect 19116 25168 19122 25220
rect 21266 25168 21272 25220
rect 21324 25168 21330 25220
rect 22278 25168 22284 25220
rect 22336 25208 22342 25220
rect 24029 25211 24087 25217
rect 24029 25208 24041 25211
rect 22336 25180 24041 25208
rect 22336 25168 22342 25180
rect 24029 25177 24041 25180
rect 24075 25177 24087 25211
rect 24029 25171 24087 25177
rect 11756 25112 12434 25140
rect 11756 25100 11762 25112
rect 15102 25100 15108 25152
rect 15160 25100 15166 25152
rect 15473 25143 15531 25149
rect 15473 25109 15485 25143
rect 15519 25140 15531 25143
rect 16666 25140 16672 25152
rect 15519 25112 16672 25140
rect 15519 25109 15531 25112
rect 15473 25103 15531 25109
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 20806 25140 20812 25152
rect 19475 25112 20812 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 20806 25100 20812 25112
rect 20864 25100 20870 25152
rect 20898 25100 20904 25152
rect 20956 25140 20962 25152
rect 21634 25140 21640 25152
rect 20956 25112 21640 25140
rect 20956 25100 20962 25112
rect 21634 25100 21640 25112
rect 21692 25140 21698 25152
rect 22097 25143 22155 25149
rect 22097 25140 22109 25143
rect 21692 25112 22109 25140
rect 21692 25100 21698 25112
rect 22097 25109 22109 25112
rect 22143 25109 22155 25143
rect 22097 25103 22155 25109
rect 22554 25100 22560 25152
rect 22612 25100 22618 25152
rect 22646 25100 22652 25152
rect 22704 25140 22710 25152
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22704 25112 22937 25140
rect 22704 25100 22710 25112
rect 22925 25109 22937 25112
rect 22971 25109 22983 25143
rect 22925 25103 22983 25109
rect 24118 25100 24124 25152
rect 24176 25140 24182 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 24176 25112 24593 25140
rect 24176 25100 24182 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 7006 24936 7012 24948
rect 6886 24908 7012 24936
rect 5994 24828 6000 24880
rect 6052 24868 6058 24880
rect 6178 24868 6184 24880
rect 6052 24840 6184 24868
rect 6052 24828 6058 24840
rect 6178 24828 6184 24840
rect 6236 24828 6242 24880
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24800 2283 24803
rect 2866 24800 2872 24812
rect 2271 24772 2872 24800
rect 2271 24769 2283 24772
rect 2225 24763 2283 24769
rect 2866 24760 2872 24772
rect 2924 24760 2930 24812
rect 6886 24800 6914 24908
rect 7006 24896 7012 24908
rect 7064 24936 7070 24948
rect 7834 24936 7840 24948
rect 7064 24908 7840 24936
rect 7064 24896 7070 24908
rect 7834 24896 7840 24908
rect 7892 24936 7898 24948
rect 7892 24908 9352 24936
rect 7892 24896 7898 24908
rect 4462 24772 6914 24800
rect 9324 24800 9352 24908
rect 10870 24896 10876 24948
rect 10928 24896 10934 24948
rect 11701 24939 11759 24945
rect 11701 24905 11713 24939
rect 11747 24905 11759 24939
rect 11701 24899 11759 24905
rect 9490 24828 9496 24880
rect 9548 24868 9554 24880
rect 10781 24871 10839 24877
rect 10781 24868 10793 24871
rect 9548 24840 10793 24868
rect 9548 24828 9554 24840
rect 10781 24837 10793 24840
rect 10827 24837 10839 24871
rect 10781 24831 10839 24837
rect 9674 24800 9680 24812
rect 9324 24786 9680 24800
rect 9338 24772 9680 24786
rect 9674 24760 9680 24772
rect 9732 24760 9738 24812
rect 9858 24760 9864 24812
rect 9916 24800 9922 24812
rect 11716 24800 11744 24899
rect 12066 24896 12072 24948
rect 12124 24896 12130 24948
rect 12434 24896 12440 24948
rect 12492 24936 12498 24948
rect 13630 24936 13636 24948
rect 12492 24908 13636 24936
rect 12492 24896 12498 24908
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 18325 24939 18383 24945
rect 18325 24905 18337 24939
rect 18371 24936 18383 24939
rect 19334 24936 19340 24948
rect 18371 24908 19340 24936
rect 18371 24905 18383 24908
rect 18325 24899 18383 24905
rect 19334 24896 19340 24908
rect 19392 24896 19398 24948
rect 19518 24896 19524 24948
rect 19576 24896 19582 24948
rect 22462 24936 22468 24948
rect 22388 24908 22468 24936
rect 9916 24772 11744 24800
rect 12161 24803 12219 24809
rect 9916 24760 9922 24772
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12526 24800 12532 24812
rect 12207 24772 12532 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12526 24760 12532 24772
rect 12584 24800 12590 24812
rect 12894 24800 12900 24812
rect 12584 24772 12900 24800
rect 12584 24760 12590 24772
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13630 24800 13636 24812
rect 13412 24772 13636 24800
rect 13412 24760 13418 24772
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 14458 24760 14464 24812
rect 14516 24800 14522 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14516 24772 14565 24800
rect 14516 24760 14522 24772
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 15930 24760 15936 24812
rect 15988 24760 15994 24812
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19613 24803 19671 24809
rect 19613 24800 19625 24803
rect 19484 24772 19625 24800
rect 19484 24760 19490 24772
rect 19613 24769 19625 24772
rect 19659 24769 19671 24803
rect 22388 24800 22416 24908
rect 22462 24896 22468 24908
rect 22520 24896 22526 24948
rect 24026 24828 24032 24880
rect 24084 24828 24090 24880
rect 19613 24763 19671 24769
rect 22296 24772 22416 24800
rect 2774 24692 2780 24744
rect 2832 24732 2838 24744
rect 3053 24735 3111 24741
rect 3053 24732 3065 24735
rect 2832 24704 3065 24732
rect 2832 24692 2838 24704
rect 3053 24701 3065 24704
rect 3099 24701 3111 24735
rect 3053 24695 3111 24701
rect 3329 24735 3387 24741
rect 3329 24701 3341 24735
rect 3375 24732 3387 24735
rect 5994 24732 6000 24744
rect 3375 24704 6000 24732
rect 3375 24701 3387 24704
rect 3329 24695 3387 24701
rect 5994 24692 6000 24704
rect 6052 24692 6058 24744
rect 6454 24692 6460 24744
rect 6512 24732 6518 24744
rect 7006 24732 7012 24744
rect 6512 24704 7012 24732
rect 6512 24692 6518 24704
rect 7006 24692 7012 24704
rect 7064 24732 7070 24744
rect 7929 24735 7987 24741
rect 7929 24732 7941 24735
rect 7064 24704 7941 24732
rect 7064 24692 7070 24704
rect 7929 24701 7941 24704
rect 7975 24701 7987 24735
rect 7929 24695 7987 24701
rect 8202 24692 8208 24744
rect 8260 24732 8266 24744
rect 10965 24735 11023 24741
rect 10965 24732 10977 24735
rect 8260 24704 10977 24732
rect 8260 24692 8266 24704
rect 10965 24701 10977 24704
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 11112 24704 12265 24732
rect 11112 24692 11118 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24732 14887 24735
rect 16206 24732 16212 24744
rect 14875 24704 16212 24732
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 16206 24692 16212 24704
rect 16264 24692 16270 24744
rect 16298 24692 16304 24744
rect 16356 24692 16362 24744
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 18417 24735 18475 24741
rect 18417 24732 18429 24735
rect 17460 24704 18429 24732
rect 17460 24692 17466 24704
rect 18417 24701 18429 24704
rect 18463 24701 18475 24735
rect 18417 24695 18475 24701
rect 18598 24692 18604 24744
rect 18656 24692 18662 24744
rect 19797 24735 19855 24741
rect 19797 24701 19809 24735
rect 19843 24732 19855 24735
rect 20622 24732 20628 24744
rect 19843 24704 20628 24732
rect 19843 24701 19855 24704
rect 19797 24695 19855 24701
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 1946 24624 1952 24676
rect 2004 24664 2010 24676
rect 2041 24667 2099 24673
rect 2041 24664 2053 24667
rect 2004 24636 2053 24664
rect 2004 24624 2010 24636
rect 2041 24633 2053 24636
rect 2087 24633 2099 24667
rect 2041 24627 2099 24633
rect 9398 24624 9404 24676
rect 9456 24664 9462 24676
rect 9677 24667 9735 24673
rect 9677 24664 9689 24667
rect 9456 24636 9689 24664
rect 9456 24624 9462 24636
rect 9677 24633 9689 24636
rect 9723 24664 9735 24667
rect 14366 24664 14372 24676
rect 9723 24636 14372 24664
rect 9723 24633 9735 24636
rect 9677 24627 9735 24633
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 22296 24664 22324 24772
rect 22462 24760 22468 24812
rect 22520 24760 22526 24812
rect 22370 24692 22376 24744
rect 22428 24732 22434 24744
rect 22557 24735 22615 24741
rect 22557 24732 22569 24735
rect 22428 24704 22569 24732
rect 22428 24692 22434 24704
rect 22557 24701 22569 24704
rect 22603 24701 22615 24735
rect 22557 24695 22615 24701
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 22756 24664 22784 24695
rect 22830 24692 22836 24744
rect 22888 24732 22894 24744
rect 23293 24735 23351 24741
rect 23293 24732 23305 24735
rect 22888 24704 23305 24732
rect 22888 24692 22894 24704
rect 23293 24701 23305 24704
rect 23339 24701 23351 24735
rect 23569 24735 23627 24741
rect 23569 24732 23581 24735
rect 23293 24695 23351 24701
rect 23400 24704 23581 24732
rect 23400 24664 23428 24704
rect 23569 24701 23581 24704
rect 23615 24732 23627 24735
rect 23658 24732 23664 24744
rect 23615 24704 23664 24732
rect 23615 24701 23627 24704
rect 23569 24695 23627 24701
rect 23658 24692 23664 24704
rect 23716 24692 23722 24744
rect 22296 24636 22416 24664
rect 22756 24636 23428 24664
rect 22388 24608 22416 24636
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 4430 24596 4436 24608
rect 4028 24568 4436 24596
rect 4028 24556 4034 24568
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 4614 24556 4620 24608
rect 4672 24596 4678 24608
rect 4801 24599 4859 24605
rect 4801 24596 4813 24599
rect 4672 24568 4813 24596
rect 4672 24556 4678 24568
rect 4801 24565 4813 24568
rect 4847 24565 4859 24599
rect 4801 24559 4859 24565
rect 7469 24599 7527 24605
rect 7469 24565 7481 24599
rect 7515 24596 7527 24599
rect 8202 24596 8208 24608
rect 7515 24568 8208 24596
rect 7515 24565 7527 24568
rect 7469 24559 7527 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 10413 24599 10471 24605
rect 10413 24565 10425 24599
rect 10459 24596 10471 24599
rect 15010 24596 15016 24608
rect 10459 24568 15016 24596
rect 10459 24565 10471 24568
rect 10413 24559 10471 24565
rect 15010 24556 15016 24568
rect 15068 24556 15074 24608
rect 17957 24599 18015 24605
rect 17957 24565 17969 24599
rect 18003 24596 18015 24599
rect 18414 24596 18420 24608
rect 18003 24568 18420 24596
rect 18003 24565 18015 24568
rect 17957 24559 18015 24565
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 19153 24599 19211 24605
rect 19153 24565 19165 24599
rect 19199 24596 19211 24599
rect 19794 24596 19800 24608
rect 19199 24568 19800 24596
rect 19199 24565 19211 24568
rect 19153 24559 19211 24565
rect 19794 24556 19800 24568
rect 19852 24556 19858 24608
rect 22094 24556 22100 24608
rect 22152 24556 22158 24608
rect 22370 24556 22376 24608
rect 22428 24596 22434 24608
rect 25041 24599 25099 24605
rect 25041 24596 25053 24599
rect 22428 24568 25053 24596
rect 22428 24556 22434 24568
rect 25041 24565 25053 24568
rect 25087 24565 25099 24599
rect 25041 24559 25099 24565
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 3145 24395 3203 24401
rect 3145 24361 3157 24395
rect 3191 24361 3203 24395
rect 3145 24355 3203 24361
rect 3160 24324 3188 24355
rect 4062 24352 4068 24404
rect 4120 24401 4126 24404
rect 4120 24395 4169 24401
rect 4120 24361 4123 24395
rect 4157 24361 4169 24395
rect 4120 24355 4169 24361
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 9490 24392 9496 24404
rect 7883 24364 9496 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 4120 24352 4126 24355
rect 9490 24352 9496 24364
rect 9548 24352 9554 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 19426 24392 19432 24404
rect 14323 24364 19432 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 22189 24395 22247 24401
rect 22189 24361 22201 24395
rect 22235 24392 22247 24395
rect 22462 24392 22468 24404
rect 22235 24364 22468 24392
rect 22235 24361 22247 24364
rect 22189 24355 22247 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 4246 24324 4252 24336
rect 3160 24296 4252 24324
rect 4246 24284 4252 24296
rect 4304 24284 4310 24336
rect 13538 24284 13544 24336
rect 13596 24324 13602 24336
rect 25133 24327 25191 24333
rect 25133 24324 25145 24327
rect 13596 24296 14872 24324
rect 13596 24284 13602 24296
rect 4430 24256 4436 24268
rect 2884 24228 4436 24256
rect 2884 24197 2912 24228
rect 4430 24216 4436 24228
rect 4488 24216 4494 24268
rect 7466 24216 7472 24268
rect 7524 24256 7530 24268
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 7524 24228 8401 24256
rect 7524 24216 7530 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 8389 24219 8447 24225
rect 9398 24216 9404 24268
rect 9456 24216 9462 24268
rect 12158 24216 12164 24268
rect 12216 24216 12222 24268
rect 12406 24228 13860 24256
rect 2869 24191 2927 24197
rect 2869 24157 2881 24191
rect 2915 24157 2927 24191
rect 4008 24191 4066 24197
rect 4008 24188 4020 24191
rect 2869 24151 2927 24157
rect 3436 24160 4020 24188
rect 2222 24080 2228 24132
rect 2280 24120 2286 24132
rect 3436 24120 3464 24160
rect 4008 24157 4020 24160
rect 4054 24157 4066 24191
rect 4008 24151 4066 24157
rect 8202 24148 8208 24200
rect 8260 24148 8266 24200
rect 9122 24148 9128 24200
rect 9180 24148 9186 24200
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12406 24188 12434 24228
rect 11931 24160 12434 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 13446 24148 13452 24200
rect 13504 24188 13510 24200
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 13504 24160 13737 24188
rect 13504 24148 13510 24160
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13832 24188 13860 24228
rect 14642 24216 14648 24268
rect 14700 24256 14706 24268
rect 14844 24265 14872 24296
rect 18248 24296 25145 24324
rect 14737 24259 14795 24265
rect 14737 24256 14749 24259
rect 14700 24228 14749 24256
rect 14700 24216 14706 24228
rect 14737 24225 14749 24228
rect 14783 24225 14795 24259
rect 14737 24219 14795 24225
rect 14829 24259 14887 24265
rect 14829 24225 14841 24259
rect 14875 24225 14887 24259
rect 14829 24219 14887 24225
rect 15746 24216 15752 24268
rect 15804 24256 15810 24268
rect 15933 24259 15991 24265
rect 15933 24256 15945 24259
rect 15804 24228 15945 24256
rect 15804 24216 15810 24228
rect 15933 24225 15945 24228
rect 15979 24225 15991 24259
rect 15933 24219 15991 24225
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 16206 24256 16212 24268
rect 16163 24228 16212 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 16206 24216 16212 24228
rect 16264 24216 16270 24268
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 18248 24265 18276 24296
rect 25133 24293 25145 24296
rect 25179 24293 25191 24327
rect 25133 24287 25191 24293
rect 18233 24259 18291 24265
rect 18233 24256 18245 24259
rect 17736 24228 18245 24256
rect 17736 24216 17742 24228
rect 18233 24225 18245 24228
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 18417 24259 18475 24265
rect 18417 24225 18429 24259
rect 18463 24256 18475 24259
rect 18506 24256 18512 24268
rect 18463 24228 18512 24256
rect 18463 24225 18475 24228
rect 18417 24219 18475 24225
rect 18506 24216 18512 24228
rect 18564 24216 18570 24268
rect 19886 24216 19892 24268
rect 19944 24216 19950 24268
rect 20073 24259 20131 24265
rect 20073 24225 20085 24259
rect 20119 24256 20131 24259
rect 20898 24256 20904 24268
rect 20119 24228 20904 24256
rect 20119 24225 20131 24228
rect 20073 24219 20131 24225
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21082 24216 21088 24268
rect 21140 24216 21146 24268
rect 21266 24216 21272 24268
rect 21324 24216 21330 24268
rect 16666 24188 16672 24200
rect 13832 24160 16672 24188
rect 13725 24151 13783 24157
rect 16666 24148 16672 24160
rect 16724 24148 16730 24200
rect 19794 24148 19800 24200
rect 19852 24148 19858 24200
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24188 22891 24191
rect 24394 24188 24400 24200
rect 22879 24160 24400 24188
rect 22879 24157 22891 24160
rect 22833 24151 22891 24157
rect 24394 24148 24400 24160
rect 24452 24148 24458 24200
rect 24762 24148 24768 24200
rect 24820 24188 24826 24200
rect 25317 24191 25375 24197
rect 25317 24188 25329 24191
rect 24820 24160 25329 24188
rect 24820 24148 24826 24160
rect 25317 24157 25329 24160
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 2280 24092 3464 24120
rect 2280 24080 2286 24092
rect 8478 24080 8484 24132
rect 8536 24120 8542 24132
rect 9490 24120 9496 24132
rect 8536 24092 9496 24120
rect 8536 24080 8542 24092
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 10410 24080 10416 24132
rect 10468 24080 10474 24132
rect 13078 24080 13084 24132
rect 13136 24120 13142 24132
rect 15841 24123 15899 24129
rect 15841 24120 15853 24123
rect 13136 24092 15853 24120
rect 13136 24080 13142 24092
rect 15841 24089 15853 24092
rect 15887 24089 15899 24123
rect 15841 24083 15899 24089
rect 18874 24080 18880 24132
rect 18932 24120 18938 24132
rect 20993 24123 21051 24129
rect 20993 24120 21005 24123
rect 18932 24092 21005 24120
rect 18932 24080 18938 24092
rect 20993 24089 21005 24092
rect 21039 24089 21051 24123
rect 20993 24083 21051 24089
rect 23845 24123 23903 24129
rect 23845 24089 23857 24123
rect 23891 24120 23903 24123
rect 24946 24120 24952 24132
rect 23891 24092 24952 24120
rect 23891 24089 23903 24092
rect 23845 24083 23903 24089
rect 24946 24080 24952 24092
rect 25004 24080 25010 24132
rect 3329 24055 3387 24061
rect 3329 24021 3341 24055
rect 3375 24052 3387 24055
rect 3418 24052 3424 24064
rect 3375 24024 3424 24052
rect 3375 24021 3387 24024
rect 3329 24015 3387 24021
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 8297 24055 8355 24061
rect 8297 24021 8309 24055
rect 8343 24052 8355 24055
rect 8386 24052 8392 24064
rect 8343 24024 8392 24052
rect 8343 24021 8355 24024
rect 8297 24015 8355 24021
rect 8386 24012 8392 24024
rect 8444 24052 8450 24064
rect 8754 24052 8760 24064
rect 8444 24024 8760 24052
rect 8444 24012 8450 24024
rect 8754 24012 8760 24024
rect 8812 24012 8818 24064
rect 10870 24012 10876 24064
rect 10928 24012 10934 24064
rect 11514 24012 11520 24064
rect 11572 24012 11578 24064
rect 11974 24012 11980 24064
rect 12032 24012 12038 24064
rect 14550 24012 14556 24064
rect 14608 24052 14614 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14608 24024 14657 24052
rect 14608 24012 14614 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 15470 24012 15476 24064
rect 15528 24012 15534 24064
rect 17770 24012 17776 24064
rect 17828 24012 17834 24064
rect 17862 24012 17868 24064
rect 17920 24052 17926 24064
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17920 24024 18153 24052
rect 17920 24012 17926 24024
rect 18141 24021 18153 24024
rect 18187 24021 18199 24055
rect 18141 24015 18199 24021
rect 18782 24012 18788 24064
rect 18840 24052 18846 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 18840 24024 19441 24052
rect 18840 24012 18846 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 20622 24012 20628 24064
rect 20680 24012 20686 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 2682 23808 2688 23860
rect 2740 23848 2746 23860
rect 4062 23848 4068 23860
rect 2740 23820 4068 23848
rect 2740 23808 2746 23820
rect 4062 23808 4068 23820
rect 4120 23848 4126 23860
rect 5534 23848 5540 23860
rect 4120 23820 5540 23848
rect 4120 23808 4126 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 5994 23808 6000 23860
rect 6052 23808 6058 23860
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 9030 23848 9036 23860
rect 8895 23820 9036 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9677 23851 9735 23857
rect 9677 23817 9689 23851
rect 9723 23848 9735 23851
rect 12253 23851 12311 23857
rect 12253 23848 12265 23851
rect 9723 23820 12265 23848
rect 9723 23817 9735 23820
rect 9677 23811 9735 23817
rect 12253 23817 12265 23820
rect 12299 23817 12311 23851
rect 12253 23811 12311 23817
rect 12342 23808 12348 23860
rect 12400 23808 12406 23860
rect 13078 23808 13084 23860
rect 13136 23808 13142 23860
rect 13446 23808 13452 23860
rect 13504 23808 13510 23860
rect 13541 23851 13599 23857
rect 13541 23817 13553 23851
rect 13587 23848 13599 23851
rect 13630 23848 13636 23860
rect 13587 23820 13636 23848
rect 13587 23817 13599 23820
rect 13541 23811 13599 23817
rect 13630 23808 13636 23820
rect 13688 23848 13694 23860
rect 14182 23848 14188 23860
rect 13688 23820 14188 23848
rect 13688 23808 13694 23820
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 23474 23848 23480 23860
rect 21140 23820 23480 23848
rect 21140 23808 21146 23820
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 2700 23780 2728 23808
rect 4982 23780 4988 23792
rect 2056 23752 2728 23780
rect 3542 23752 4988 23780
rect 2056 23721 2084 23752
rect 4982 23740 4988 23752
rect 5040 23740 5046 23792
rect 6638 23740 6644 23792
rect 6696 23780 6702 23792
rect 11606 23780 11612 23792
rect 6696 23752 11612 23780
rect 6696 23740 6702 23752
rect 11606 23740 11612 23752
rect 11664 23780 11670 23792
rect 11974 23780 11980 23792
rect 11664 23752 11980 23780
rect 11664 23740 11670 23752
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 24854 23780 24860 23792
rect 22296 23752 24860 23780
rect 2041 23715 2099 23721
rect 2041 23681 2053 23715
rect 2087 23681 2099 23715
rect 2041 23675 2099 23681
rect 4062 23672 4068 23724
rect 4120 23712 4126 23724
rect 4249 23715 4307 23721
rect 4249 23712 4261 23715
rect 4120 23684 4261 23712
rect 4120 23672 4126 23684
rect 4249 23681 4261 23684
rect 4295 23681 4307 23715
rect 7098 23712 7104 23724
rect 4249 23675 4307 23681
rect 5552 23684 7104 23712
rect 2317 23647 2375 23653
rect 2317 23613 2329 23647
rect 2363 23644 2375 23647
rect 4614 23644 4620 23656
rect 2363 23616 4620 23644
rect 2363 23613 2375 23616
rect 2317 23607 2375 23613
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 4982 23604 4988 23656
rect 5040 23644 5046 23656
rect 5552 23644 5580 23684
rect 7098 23672 7104 23684
rect 7156 23672 7162 23724
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23712 8999 23715
rect 10045 23715 10103 23721
rect 8987 23684 9352 23712
rect 8987 23681 8999 23684
rect 8941 23675 8999 23681
rect 5040 23616 5580 23644
rect 5040 23604 5046 23616
rect 9030 23604 9036 23656
rect 9088 23604 9094 23656
rect 3789 23511 3847 23517
rect 3789 23477 3801 23511
rect 3835 23508 3847 23511
rect 4246 23508 4252 23520
rect 3835 23480 4252 23508
rect 3835 23477 3847 23480
rect 3789 23471 3847 23477
rect 4246 23468 4252 23480
rect 4304 23468 4310 23520
rect 4512 23511 4570 23517
rect 4512 23477 4524 23511
rect 4558 23508 4570 23511
rect 5810 23508 5816 23520
rect 4558 23480 5816 23508
rect 4558 23477 4570 23480
rect 4512 23471 4570 23477
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 8478 23468 8484 23520
rect 8536 23468 8542 23520
rect 9324 23508 9352 23684
rect 10045 23681 10057 23715
rect 10091 23712 10103 23715
rect 11057 23715 11115 23721
rect 11057 23712 11069 23715
rect 10091 23684 11069 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 11057 23681 11069 23684
rect 11103 23681 11115 23715
rect 11057 23675 11115 23681
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 16482 23712 16488 23724
rect 13596 23684 16488 23712
rect 13596 23672 13602 23684
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 22296 23721 22324 23752
rect 24854 23740 24860 23752
rect 24912 23740 24918 23792
rect 25130 23740 25136 23792
rect 25188 23740 25194 23792
rect 22281 23715 22339 23721
rect 22281 23681 22293 23715
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 24118 23672 24124 23724
rect 24176 23672 24182 23724
rect 9490 23604 9496 23656
rect 9548 23644 9554 23656
rect 10137 23647 10195 23653
rect 10137 23644 10149 23647
rect 9548 23616 10149 23644
rect 9548 23604 9554 23616
rect 10137 23613 10149 23616
rect 10183 23613 10195 23647
rect 10137 23607 10195 23613
rect 10229 23647 10287 23653
rect 10229 23613 10241 23647
rect 10275 23613 10287 23647
rect 10229 23607 10287 23613
rect 9398 23536 9404 23588
rect 9456 23576 9462 23588
rect 10244 23576 10272 23607
rect 10870 23604 10876 23656
rect 10928 23644 10934 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 10928 23616 12449 23644
rect 10928 23604 10934 23616
rect 12437 23613 12449 23616
rect 12483 23613 12495 23647
rect 12437 23607 12495 23613
rect 13725 23647 13783 23653
rect 13725 23613 13737 23647
rect 13771 23644 13783 23647
rect 16390 23644 16396 23656
rect 13771 23616 16396 23644
rect 13771 23613 13783 23616
rect 13725 23607 13783 23613
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 23293 23647 23351 23653
rect 23293 23613 23305 23647
rect 23339 23644 23351 23647
rect 23382 23644 23388 23656
rect 23339 23616 23388 23644
rect 23339 23613 23351 23616
rect 23293 23607 23351 23613
rect 23382 23604 23388 23616
rect 23440 23604 23446 23656
rect 11974 23576 11980 23588
rect 9456 23548 10272 23576
rect 10336 23548 11980 23576
rect 9456 23536 9462 23548
rect 10336 23508 10364 23548
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 9324 23480 10364 23508
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 15286 23508 15292 23520
rect 11931 23480 15292 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 3326 23264 3332 23316
rect 3384 23304 3390 23316
rect 4065 23307 4123 23313
rect 4065 23304 4077 23307
rect 3384 23276 4077 23304
rect 3384 23264 3390 23276
rect 4065 23273 4077 23276
rect 4111 23273 4123 23307
rect 4065 23267 4123 23273
rect 5810 23264 5816 23316
rect 5868 23304 5874 23316
rect 6822 23304 6828 23316
rect 5868 23276 6828 23304
rect 5868 23264 5874 23276
rect 6822 23264 6828 23276
rect 6880 23304 6886 23316
rect 7285 23307 7343 23313
rect 7285 23304 7297 23307
rect 6880 23276 7297 23304
rect 6880 23264 6886 23276
rect 7285 23273 7297 23276
rect 7331 23273 7343 23307
rect 18874 23304 18880 23316
rect 7285 23267 7343 23273
rect 17420 23276 18880 23304
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 16206 23236 16212 23248
rect 15703 23208 16212 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 16206 23196 16212 23208
rect 16264 23196 16270 23248
rect 1302 23128 1308 23180
rect 1360 23168 1366 23180
rect 2041 23171 2099 23177
rect 2041 23168 2053 23171
rect 1360 23140 2053 23168
rect 1360 23128 1366 23140
rect 2041 23137 2053 23140
rect 2087 23137 2099 23171
rect 2041 23131 2099 23137
rect 5534 23128 5540 23180
rect 5592 23168 5598 23180
rect 7006 23168 7012 23180
rect 5592 23140 7012 23168
rect 5592 23128 5598 23140
rect 7006 23128 7012 23140
rect 7064 23168 7070 23180
rect 7834 23168 7840 23180
rect 7064 23140 7840 23168
rect 7064 23128 7070 23140
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 10134 23128 10140 23180
rect 10192 23128 10198 23180
rect 16298 23128 16304 23180
rect 16356 23128 16362 23180
rect 17420 23177 17448 23276
rect 18874 23264 18880 23276
rect 18932 23264 18938 23316
rect 19518 23264 19524 23316
rect 19576 23304 19582 23316
rect 20714 23304 20720 23316
rect 19576 23276 20720 23304
rect 19576 23264 19582 23276
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 20993 23239 21051 23245
rect 20993 23205 21005 23239
rect 21039 23236 21051 23239
rect 22738 23236 22744 23248
rect 21039 23208 22744 23236
rect 21039 23205 21051 23208
rect 20993 23199 21051 23205
rect 22738 23196 22744 23208
rect 22796 23196 22802 23248
rect 17405 23171 17463 23177
rect 17405 23137 17417 23171
rect 17451 23137 17463 23171
rect 17405 23131 17463 23137
rect 17589 23171 17647 23177
rect 17589 23137 17601 23171
rect 17635 23168 17647 23171
rect 18506 23168 18512 23180
rect 17635 23140 18512 23168
rect 17635 23137 17647 23140
rect 17589 23131 17647 23137
rect 18506 23128 18512 23140
rect 18564 23168 18570 23180
rect 18874 23168 18880 23180
rect 18564 23140 18880 23168
rect 18564 23128 18570 23140
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 21910 23128 21916 23180
rect 21968 23128 21974 23180
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 22370 23168 22376 23180
rect 22051 23140 22376 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 2682 23100 2688 23112
rect 1811 23072 2688 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23100 9919 23103
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 9907 23072 10885 23100
rect 9907 23069 9919 23072
rect 9861 23063 9919 23069
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 4264 23032 4292 23063
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15528 23072 16037 23100
rect 15528 23060 15534 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 16117 23103 16175 23109
rect 16117 23069 16129 23103
rect 16163 23100 16175 23103
rect 16574 23100 16580 23112
rect 16163 23072 16580 23100
rect 16163 23069 16175 23072
rect 16117 23063 16175 23069
rect 16574 23060 16580 23072
rect 16632 23060 16638 23112
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23100 21879 23103
rect 22094 23100 22100 23112
rect 21867 23072 22100 23100
rect 21867 23069 21879 23072
rect 21821 23063 21879 23069
rect 5718 23032 5724 23044
rect 4264 23004 5724 23032
rect 5718 22992 5724 23004
rect 5776 22992 5782 23044
rect 5813 23035 5871 23041
rect 5813 23001 5825 23035
rect 5859 23001 5871 23035
rect 7098 23032 7104 23044
rect 7038 23004 7104 23032
rect 5813 22995 5871 23001
rect 5828 22964 5856 22995
rect 7098 22992 7104 23004
rect 7156 23032 7162 23044
rect 9674 23032 9680 23044
rect 7156 23004 9680 23032
rect 7156 22992 7162 23004
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 13722 22992 13728 23044
rect 13780 23032 13786 23044
rect 18340 23032 18368 23063
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23566 23100 23572 23112
rect 22879 23072 23572 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 23566 23060 23572 23072
rect 23624 23060 23630 23112
rect 13780 23004 18368 23032
rect 23845 23035 23903 23041
rect 13780 22992 13786 23004
rect 23845 23001 23857 23035
rect 23891 23032 23903 23035
rect 26050 23032 26056 23044
rect 23891 23004 26056 23032
rect 23891 23001 23903 23004
rect 23845 22995 23903 23001
rect 26050 22992 26056 23004
rect 26108 22992 26114 23044
rect 8294 22964 8300 22976
rect 5828 22936 8300 22964
rect 8294 22924 8300 22936
rect 8352 22964 8358 22976
rect 9030 22964 9036 22976
rect 8352 22936 9036 22964
rect 8352 22924 8358 22936
rect 9030 22924 9036 22936
rect 9088 22924 9094 22976
rect 9490 22924 9496 22976
rect 9548 22924 9554 22976
rect 9953 22967 10011 22973
rect 9953 22933 9965 22967
rect 9999 22964 10011 22967
rect 11422 22964 11428 22976
rect 9999 22936 11428 22964
rect 9999 22933 10011 22936
rect 9953 22927 10011 22933
rect 11422 22924 11428 22936
rect 11480 22964 11486 22976
rect 12250 22964 12256 22976
rect 11480 22936 12256 22964
rect 11480 22924 11486 22936
rect 12250 22924 12256 22936
rect 12308 22924 12314 22976
rect 14458 22924 14464 22976
rect 14516 22964 14522 22976
rect 16758 22964 16764 22976
rect 14516 22936 16764 22964
rect 14516 22924 14522 22936
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 16945 22967 17003 22973
rect 16945 22933 16957 22967
rect 16991 22964 17003 22967
rect 17218 22964 17224 22976
rect 16991 22936 17224 22964
rect 16991 22933 17003 22936
rect 16945 22927 17003 22933
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 17310 22924 17316 22976
rect 17368 22924 17374 22976
rect 18141 22967 18199 22973
rect 18141 22933 18153 22967
rect 18187 22964 18199 22967
rect 19242 22964 19248 22976
rect 18187 22936 19248 22964
rect 18187 22933 18199 22936
rect 18141 22927 18199 22933
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21453 22967 21511 22973
rect 21453 22964 21465 22967
rect 21232 22936 21465 22964
rect 21232 22924 21238 22936
rect 21453 22933 21465 22936
rect 21499 22933 21511 22967
rect 21453 22927 21511 22933
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22646 22964 22652 22976
rect 22152 22936 22652 22964
rect 22152 22924 22158 22936
rect 22646 22924 22652 22936
rect 22704 22924 22710 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 1949 22763 2007 22769
rect 1949 22760 1961 22763
rect 1820 22732 1961 22760
rect 1820 22720 1826 22732
rect 1949 22729 1961 22732
rect 1995 22729 2007 22763
rect 1949 22723 2007 22729
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 3237 22763 3295 22769
rect 3237 22760 3249 22763
rect 2924 22732 3249 22760
rect 2924 22720 2930 22732
rect 3237 22729 3249 22732
rect 3283 22729 3295 22763
rect 3237 22723 3295 22729
rect 3878 22720 3884 22772
rect 3936 22760 3942 22772
rect 4019 22763 4077 22769
rect 4019 22760 4031 22763
rect 3936 22732 4031 22760
rect 3936 22720 3942 22732
rect 4019 22729 4031 22732
rect 4065 22729 4077 22763
rect 10042 22760 10048 22772
rect 4019 22723 4077 22729
rect 7484 22732 10048 22760
rect 7484 22701 7512 22732
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 12529 22763 12587 22769
rect 12529 22729 12541 22763
rect 12575 22760 12587 22763
rect 14458 22760 14464 22772
rect 12575 22732 14464 22760
rect 12575 22729 12587 22732
rect 12529 22723 12587 22729
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 14550 22720 14556 22772
rect 14608 22760 14614 22772
rect 15105 22763 15163 22769
rect 15105 22760 15117 22763
rect 14608 22732 15117 22760
rect 14608 22720 14614 22732
rect 15105 22729 15117 22732
rect 15151 22760 15163 22763
rect 15654 22760 15660 22772
rect 15151 22732 15660 22760
rect 15151 22729 15163 22732
rect 15105 22723 15163 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16448 22732 18460 22760
rect 16448 22720 16454 22732
rect 7469 22695 7527 22701
rect 7469 22661 7481 22695
rect 7515 22661 7527 22695
rect 7469 22655 7527 22661
rect 9674 22652 9680 22704
rect 9732 22652 9738 22704
rect 12618 22652 12624 22704
rect 12676 22692 12682 22704
rect 13630 22692 13636 22704
rect 12676 22664 13636 22692
rect 12676 22652 12682 22664
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 15930 22692 15936 22704
rect 14858 22664 15936 22692
rect 15930 22652 15936 22664
rect 15988 22692 15994 22704
rect 16482 22692 16488 22704
rect 15988 22664 16488 22692
rect 15988 22652 15994 22664
rect 16482 22652 16488 22664
rect 16540 22692 16546 22704
rect 18432 22692 18460 22732
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 18564 22732 18613 22760
rect 18564 22720 18570 22732
rect 18601 22729 18613 22732
rect 18647 22729 18659 22763
rect 18601 22723 18659 22729
rect 18708 22732 21128 22760
rect 18708 22692 18736 22732
rect 16540 22664 17618 22692
rect 18432 22664 18736 22692
rect 16540 22652 16546 22664
rect 19058 22652 19064 22704
rect 19116 22692 19122 22704
rect 19794 22692 19800 22704
rect 19116 22664 19800 22692
rect 19116 22652 19122 22664
rect 19794 22652 19800 22664
rect 19852 22652 19858 22704
rect 21100 22701 21128 22732
rect 22370 22720 22376 22772
rect 22428 22720 22434 22772
rect 23474 22720 23480 22772
rect 23532 22760 23538 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 23532 22732 24777 22760
rect 23532 22720 23538 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 21085 22695 21143 22701
rect 21085 22661 21097 22695
rect 21131 22661 21143 22695
rect 22388 22692 22416 22720
rect 23293 22695 23351 22701
rect 23293 22692 23305 22695
rect 21085 22655 21143 22661
rect 22066 22664 23305 22692
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22624 2191 22627
rect 2866 22624 2872 22636
rect 2179 22596 2872 22624
rect 2179 22593 2191 22596
rect 2133 22587 2191 22593
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3916 22627 3974 22633
rect 3916 22624 3928 22627
rect 3568 22596 3928 22624
rect 3568 22584 3574 22596
rect 3916 22593 3928 22596
rect 3962 22593 3974 22627
rect 3916 22587 3974 22593
rect 5626 22584 5632 22636
rect 5684 22584 5690 22636
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22624 5779 22627
rect 7650 22624 7656 22636
rect 5767 22596 7656 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 12894 22624 12900 22636
rect 12636 22596 12900 22624
rect 2593 22559 2651 22565
rect 2593 22525 2605 22559
rect 2639 22525 2651 22559
rect 2593 22519 2651 22525
rect 2608 22488 2636 22519
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 3418 22556 3424 22568
rect 2832 22528 3424 22556
rect 2832 22516 2838 22528
rect 3418 22516 3424 22528
rect 3476 22516 3482 22568
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 5994 22556 6000 22568
rect 5951 22528 6000 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7834 22516 7840 22568
rect 7892 22556 7898 22568
rect 8205 22559 8263 22565
rect 8205 22556 8217 22559
rect 7892 22528 8217 22556
rect 7892 22516 7898 22528
rect 8205 22525 8217 22528
rect 8251 22525 8263 22559
rect 8205 22519 8263 22525
rect 8849 22559 8907 22565
rect 8849 22525 8861 22559
rect 8895 22556 8907 22559
rect 9125 22559 9183 22565
rect 8895 22528 8984 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 4798 22488 4804 22500
rect 2608 22460 4804 22488
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 5261 22423 5319 22429
rect 5261 22420 5273 22423
rect 4212 22392 5273 22420
rect 4212 22380 4218 22392
rect 5261 22389 5273 22392
rect 5307 22389 5319 22423
rect 8956 22420 8984 22528
rect 9125 22525 9137 22559
rect 9171 22556 9183 22559
rect 10870 22556 10876 22568
rect 9171 22528 10876 22556
rect 9171 22525 9183 22528
rect 9125 22519 9183 22525
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 11790 22516 11796 22568
rect 11848 22556 11854 22568
rect 12636 22565 12664 22596
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 15749 22627 15807 22633
rect 15749 22593 15761 22627
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 12621 22559 12679 22565
rect 11848 22528 12388 22556
rect 11848 22516 11854 22528
rect 11808 22488 11836 22516
rect 10152 22460 11836 22488
rect 9122 22420 9128 22432
rect 8956 22392 9128 22420
rect 5261 22383 5319 22389
rect 9122 22380 9128 22392
rect 9180 22420 9186 22432
rect 10152 22420 10180 22460
rect 12066 22448 12072 22500
rect 12124 22488 12130 22500
rect 12360 22488 12388 22528
rect 12621 22525 12633 22559
rect 12667 22525 12679 22559
rect 12621 22519 12679 22525
rect 12802 22516 12808 22568
rect 12860 22516 12866 22568
rect 13354 22516 13360 22568
rect 13412 22516 13418 22568
rect 15764 22556 15792 22587
rect 16850 22584 16856 22636
rect 16908 22584 16914 22636
rect 14660 22528 15792 22556
rect 13372 22488 13400 22516
rect 12124 22460 12296 22488
rect 12360 22460 13400 22488
rect 12124 22448 12130 22460
rect 9180 22392 10180 22420
rect 9180 22380 9186 22392
rect 10594 22380 10600 22432
rect 10652 22420 10658 22432
rect 10962 22420 10968 22432
rect 10652 22392 10968 22420
rect 10652 22380 10658 22392
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 12158 22380 12164 22432
rect 12216 22380 12222 22432
rect 12268 22420 12296 22460
rect 14660 22420 14688 22528
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17586 22556 17592 22568
rect 16816 22528 17592 22556
rect 16816 22516 16822 22528
rect 17586 22516 17592 22528
rect 17644 22516 17650 22568
rect 18966 22516 18972 22568
rect 19024 22556 19030 22568
rect 19061 22559 19119 22565
rect 19061 22556 19073 22559
rect 19024 22528 19073 22556
rect 19024 22516 19030 22528
rect 19061 22525 19073 22528
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 19334 22516 19340 22568
rect 19392 22516 19398 22568
rect 21266 22516 21272 22568
rect 21324 22556 21330 22568
rect 22066 22556 22094 22664
rect 23293 22661 23305 22664
rect 23339 22661 23351 22695
rect 23293 22655 23351 22661
rect 24026 22652 24032 22704
rect 24084 22652 24090 22704
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 22244 22596 22385 22624
rect 22244 22584 22250 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 21324 22528 22094 22556
rect 21324 22516 21330 22528
rect 22646 22516 22652 22568
rect 22704 22556 22710 22568
rect 22830 22556 22836 22568
rect 22704 22528 22836 22556
rect 22704 22516 22710 22528
rect 22830 22516 22836 22528
rect 22888 22556 22894 22568
rect 23017 22559 23075 22565
rect 23017 22556 23029 22559
rect 22888 22528 23029 22556
rect 22888 22516 22894 22528
rect 23017 22525 23029 22528
rect 23063 22525 23075 22559
rect 23017 22519 23075 22525
rect 12268 22392 14688 22420
rect 15565 22423 15623 22429
rect 15565 22389 15577 22423
rect 15611 22420 15623 22423
rect 15930 22420 15936 22432
rect 15611 22392 15936 22420
rect 15611 22389 15623 22392
rect 15565 22383 15623 22389
rect 15930 22380 15936 22392
rect 15988 22380 15994 22432
rect 17126 22429 17132 22432
rect 17116 22423 17132 22429
rect 17116 22389 17128 22423
rect 17184 22420 17190 22432
rect 17678 22420 17684 22432
rect 17184 22392 17684 22420
rect 17116 22383 17132 22389
rect 17126 22380 17132 22383
rect 17184 22380 17190 22392
rect 17678 22380 17684 22392
rect 17736 22380 17742 22432
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19058 22420 19064 22432
rect 18932 22392 19064 22420
rect 18932 22380 18938 22392
rect 19058 22380 19064 22392
rect 19116 22380 19122 22432
rect 19794 22380 19800 22432
rect 19852 22420 19858 22432
rect 20346 22420 20352 22432
rect 19852 22392 20352 22420
rect 19852 22380 19858 22392
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 22462 22380 22468 22432
rect 22520 22380 22526 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 2682 22176 2688 22228
rect 2740 22176 2746 22228
rect 5626 22176 5632 22228
rect 5684 22216 5690 22228
rect 6089 22219 6147 22225
rect 6089 22216 6101 22219
rect 5684 22188 6101 22216
rect 5684 22176 5690 22188
rect 6089 22185 6101 22188
rect 6135 22185 6147 22219
rect 6089 22179 6147 22185
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7524 22188 7788 22216
rect 7524 22176 7530 22188
rect 6822 22148 6828 22160
rect 6748 22120 6828 22148
rect 3602 22080 3608 22092
rect 2240 22052 3608 22080
rect 2240 22021 2268 22052
rect 3602 22040 3608 22052
rect 3660 22040 3666 22092
rect 6748 22089 6776 22120
rect 6822 22108 6828 22120
rect 6880 22148 6886 22160
rect 7558 22148 7564 22160
rect 6880 22120 7564 22148
rect 6880 22108 6886 22120
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 7760 22148 7788 22188
rect 8938 22176 8944 22228
rect 8996 22216 9002 22228
rect 10226 22216 10232 22228
rect 8996 22188 10232 22216
rect 8996 22176 9002 22188
rect 10226 22176 10232 22188
rect 10284 22216 10290 22228
rect 18966 22216 18972 22228
rect 10284 22188 12388 22216
rect 10284 22176 10290 22188
rect 7760 22120 7880 22148
rect 6733 22083 6791 22089
rect 6733 22049 6745 22083
rect 6779 22080 6791 22083
rect 6779 22052 6813 22080
rect 6779 22049 6791 22052
rect 6733 22043 6791 22049
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7374 22080 7380 22092
rect 7156 22052 7380 22080
rect 7156 22040 7162 22052
rect 7374 22040 7380 22052
rect 7432 22040 7438 22092
rect 7466 22040 7472 22092
rect 7524 22040 7530 22092
rect 7852 22089 7880 22120
rect 11606 22108 11612 22160
rect 11664 22148 11670 22160
rect 11664 22120 12296 22148
rect 11664 22108 11670 22120
rect 7837 22083 7895 22089
rect 7837 22049 7849 22083
rect 7883 22080 7895 22083
rect 11425 22083 11483 22089
rect 7883 22052 7917 22080
rect 7883 22049 7895 22052
rect 7837 22043 7895 22049
rect 11425 22049 11437 22083
rect 11471 22080 11483 22083
rect 11790 22080 11796 22092
rect 11471 22052 11796 22080
rect 11471 22049 11483 22052
rect 11425 22043 11483 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 2866 21972 2872 22024
rect 2924 21972 2930 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7484 22012 7512 22040
rect 7064 21984 7512 22012
rect 7653 22015 7711 22021
rect 7064 21972 7070 21984
rect 7653 21981 7665 22015
rect 7699 22012 7711 22015
rect 9490 22012 9496 22024
rect 7699 21984 9496 22012
rect 7699 21981 7711 21984
rect 7653 21975 7711 21981
rect 9490 21972 9496 21984
rect 9548 21972 9554 22024
rect 12268 22012 12296 22120
rect 12360 22080 12388 22188
rect 12544 22188 14872 22216
rect 12544 22089 12572 22188
rect 14274 22108 14280 22160
rect 14332 22108 14338 22160
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 12360 22052 12449 22080
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 12529 22083 12587 22089
rect 12529 22049 12541 22083
rect 12575 22049 12587 22083
rect 13630 22080 13636 22092
rect 12529 22043 12587 22049
rect 13280 22052 13636 22080
rect 12544 22012 12572 22043
rect 12268 21984 12572 22012
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 13280 22012 13308 22052
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 14844 22089 14872 22188
rect 16960 22188 18972 22216
rect 16960 22092 16988 22188
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 20422 22219 20480 22225
rect 20422 22216 20434 22219
rect 19116 22188 20434 22216
rect 19116 22176 19122 22188
rect 20422 22185 20434 22188
rect 20468 22216 20480 22219
rect 22922 22216 22928 22228
rect 20468 22188 22928 22216
rect 20468 22185 20480 22188
rect 20422 22179 20480 22185
rect 22922 22176 22928 22188
rect 22980 22176 22986 22228
rect 17405 22151 17463 22157
rect 17405 22117 17417 22151
rect 17451 22148 17463 22151
rect 17678 22148 17684 22160
rect 17451 22120 17684 22148
rect 17451 22117 17463 22120
rect 17405 22111 17463 22117
rect 17678 22108 17684 22120
rect 17736 22108 17742 22160
rect 19702 22148 19708 22160
rect 18800 22120 19708 22148
rect 14829 22083 14887 22089
rect 14829 22049 14841 22083
rect 14875 22080 14887 22083
rect 15657 22083 15715 22089
rect 14875 22052 14909 22080
rect 14875 22049 14887 22052
rect 14829 22043 14887 22049
rect 15657 22049 15669 22083
rect 15703 22080 15715 22083
rect 16942 22080 16948 22092
rect 15703 22052 16948 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 16942 22040 16948 22052
rect 17000 22040 17006 22092
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 18800 22089 18828 22120
rect 19702 22108 19708 22120
rect 19760 22148 19766 22160
rect 20070 22148 20076 22160
rect 19760 22120 20076 22148
rect 19760 22108 19766 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 22646 22108 22652 22160
rect 22704 22108 22710 22160
rect 18601 22083 18659 22089
rect 18601 22080 18613 22083
rect 17828 22052 18613 22080
rect 17828 22040 17834 22052
rect 18601 22049 18613 22052
rect 18647 22049 18659 22083
rect 18601 22043 18659 22049
rect 18785 22083 18843 22089
rect 18785 22049 18797 22083
rect 18831 22080 18843 22083
rect 18831 22052 18865 22080
rect 18831 22049 18843 22052
rect 18785 22043 18843 22049
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 20165 22083 20223 22089
rect 20165 22080 20177 22083
rect 19668 22052 20177 22080
rect 19668 22040 19674 22052
rect 20165 22049 20177 22052
rect 20211 22080 20223 22083
rect 22664 22080 22692 22108
rect 20211 22052 22692 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 12676 21984 13308 22012
rect 13357 22015 13415 22021
rect 12676 21972 12682 21984
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 13906 22012 13912 22024
rect 13403 21984 13912 22012
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14645 22015 14703 22021
rect 14645 21981 14657 22015
rect 14691 22012 14703 22015
rect 15194 22012 15200 22024
rect 14691 21984 15200 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 18509 22015 18567 22021
rect 18509 22012 18521 22015
rect 17276 21984 18521 22012
rect 17276 21972 17282 21984
rect 18509 21981 18521 21984
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 22012 22891 22015
rect 24210 22012 24216 22024
rect 22879 21984 24216 22012
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 24210 21972 24216 21984
rect 24268 21972 24274 22024
rect 6457 21947 6515 21953
rect 6457 21913 6469 21947
rect 6503 21944 6515 21947
rect 8478 21944 8484 21956
rect 6503 21916 8484 21944
rect 6503 21913 6515 21916
rect 6457 21907 6515 21913
rect 8478 21904 8484 21916
rect 8536 21904 8542 21956
rect 10042 21904 10048 21956
rect 10100 21944 10106 21956
rect 10597 21947 10655 21953
rect 10597 21944 10609 21947
rect 10100 21916 10609 21944
rect 10100 21904 10106 21916
rect 10597 21913 10609 21916
rect 10643 21944 10655 21947
rect 15838 21944 15844 21956
rect 10643 21916 15844 21944
rect 10643 21913 10655 21916
rect 10597 21907 10655 21913
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 15933 21947 15991 21953
rect 15933 21913 15945 21947
rect 15979 21944 15991 21947
rect 16022 21944 16028 21956
rect 15979 21916 16028 21944
rect 15979 21913 15991 21916
rect 15933 21907 15991 21913
rect 16022 21904 16028 21916
rect 16080 21904 16086 21956
rect 16482 21904 16488 21956
rect 16540 21904 16546 21956
rect 20346 21904 20352 21956
rect 20404 21944 20410 21956
rect 23845 21947 23903 21953
rect 20404 21916 20930 21944
rect 20404 21904 20410 21916
rect 23845 21913 23857 21947
rect 23891 21944 23903 21947
rect 24946 21944 24952 21956
rect 23891 21916 24952 21944
rect 23891 21913 23903 21916
rect 23845 21907 23903 21913
rect 24946 21904 24952 21916
rect 25004 21904 25010 21956
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 2041 21879 2099 21885
rect 2041 21876 2053 21879
rect 1820 21848 2053 21876
rect 1820 21836 1826 21848
rect 2041 21845 2053 21848
rect 2087 21845 2099 21879
rect 2041 21839 2099 21845
rect 6546 21836 6552 21888
rect 6604 21836 6610 21888
rect 7282 21836 7288 21888
rect 7340 21836 7346 21888
rect 7742 21836 7748 21888
rect 7800 21836 7806 21888
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 11977 21879 12035 21885
rect 11977 21876 11989 21879
rect 9548 21848 11989 21876
rect 9548 21836 9554 21848
rect 11977 21845 11989 21848
rect 12023 21845 12035 21879
rect 11977 21839 12035 21845
rect 12342 21836 12348 21888
rect 12400 21836 12406 21888
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 13173 21879 13231 21885
rect 13173 21876 13185 21879
rect 12768 21848 13185 21876
rect 12768 21836 12774 21848
rect 13173 21845 13185 21848
rect 13219 21845 13231 21879
rect 13173 21839 13231 21845
rect 13262 21836 13268 21888
rect 13320 21876 13326 21888
rect 14642 21876 14648 21888
rect 13320 21848 14648 21876
rect 13320 21836 13326 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14734 21836 14740 21888
rect 14792 21836 14798 21888
rect 14826 21836 14832 21888
rect 14884 21876 14890 21888
rect 16114 21876 16120 21888
rect 14884 21848 16120 21876
rect 14884 21836 14890 21848
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 18141 21879 18199 21885
rect 18141 21876 18153 21879
rect 17920 21848 18153 21876
rect 17920 21836 17926 21848
rect 18141 21845 18153 21848
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 20162 21876 20168 21888
rect 19944 21848 20168 21876
rect 19944 21836 19950 21848
rect 20162 21836 20168 21848
rect 20220 21876 20226 21888
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 20220 21848 21925 21876
rect 20220 21836 20226 21848
rect 21913 21845 21925 21848
rect 21959 21845 21971 21879
rect 21913 21839 21971 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2958 21632 2964 21684
rect 3016 21672 3022 21684
rect 3145 21675 3203 21681
rect 3145 21672 3157 21675
rect 3016 21644 3157 21672
rect 3016 21632 3022 21644
rect 3145 21641 3157 21644
rect 3191 21641 3203 21675
rect 3145 21635 3203 21641
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 6549 21675 6607 21681
rect 6549 21672 6561 21675
rect 5776 21644 6561 21672
rect 5776 21632 5782 21644
rect 6549 21641 6561 21644
rect 6595 21641 6607 21675
rect 6549 21635 6607 21641
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7282 21672 7288 21684
rect 6963 21644 7288 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 7745 21675 7803 21681
rect 7745 21672 7757 21675
rect 7708 21644 7757 21672
rect 7708 21632 7714 21644
rect 7745 21641 7757 21644
rect 7791 21641 7803 21675
rect 7745 21635 7803 21641
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 14734 21672 14740 21684
rect 10744 21644 14740 21672
rect 10744 21632 10750 21644
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 17494 21672 17500 21684
rect 15252 21644 17500 21672
rect 15252 21632 15258 21644
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 19334 21632 19340 21684
rect 19392 21672 19398 21684
rect 21361 21675 21419 21681
rect 21361 21672 21373 21675
rect 19392 21644 21373 21672
rect 19392 21632 19398 21644
rect 21361 21641 21373 21644
rect 21407 21641 21419 21675
rect 23750 21672 23756 21684
rect 21361 21635 21419 21641
rect 22066 21644 23152 21672
rect 2774 21564 2780 21616
rect 2832 21604 2838 21616
rect 3326 21604 3332 21616
rect 2832 21576 3332 21604
rect 2832 21564 2838 21576
rect 3326 21564 3332 21576
rect 3384 21564 3390 21616
rect 7009 21607 7067 21613
rect 7009 21573 7021 21607
rect 7055 21604 7067 21607
rect 9122 21604 9128 21616
rect 7055 21576 9128 21604
rect 7055 21573 7067 21576
rect 7009 21567 7067 21573
rect 9122 21564 9128 21576
rect 9180 21564 9186 21616
rect 10321 21607 10379 21613
rect 10321 21573 10333 21607
rect 10367 21604 10379 21607
rect 13262 21604 13268 21616
rect 10367 21576 13268 21604
rect 10367 21573 10379 21576
rect 10321 21567 10379 21573
rect 13262 21564 13268 21576
rect 13320 21564 13326 21616
rect 13906 21564 13912 21616
rect 13964 21604 13970 21616
rect 14369 21607 14427 21613
rect 14369 21604 14381 21607
rect 13964 21576 14381 21604
rect 13964 21564 13970 21576
rect 14369 21573 14381 21576
rect 14415 21573 14427 21607
rect 14369 21567 14427 21573
rect 15838 21564 15844 21616
rect 15896 21604 15902 21616
rect 18141 21607 18199 21613
rect 18141 21604 18153 21607
rect 15896 21576 18153 21604
rect 15896 21564 15902 21576
rect 18141 21573 18153 21576
rect 18187 21604 18199 21607
rect 18322 21604 18328 21616
rect 18187 21576 18328 21604
rect 18187 21573 18199 21576
rect 18141 21567 18199 21573
rect 18322 21564 18328 21576
rect 18380 21564 18386 21616
rect 18966 21564 18972 21616
rect 19024 21564 19030 21616
rect 19886 21564 19892 21616
rect 19944 21564 19950 21616
rect 20346 21564 20352 21616
rect 20404 21564 20410 21616
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 3786 21536 3792 21548
rect 2547 21508 3792 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 3786 21496 3792 21508
rect 3844 21496 3850 21548
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 4154 21536 4160 21548
rect 3927 21508 4160 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4430 21496 4436 21548
rect 4488 21496 4494 21548
rect 8110 21496 8116 21548
rect 8168 21496 8174 21548
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21536 8263 21539
rect 10226 21536 10232 21548
rect 8251 21508 10232 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 11698 21536 11704 21548
rect 10428 21508 11704 21536
rect 10428 21480 10456 21508
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 12342 21496 12348 21548
rect 12400 21536 12406 21548
rect 12894 21536 12900 21548
rect 12400 21508 12900 21536
rect 12400 21496 12406 21508
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21536 13139 21539
rect 13722 21536 13728 21548
rect 13127 21508 13728 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 2222 21428 2228 21480
rect 2280 21468 2286 21480
rect 2685 21471 2743 21477
rect 2685 21468 2697 21471
rect 2280 21440 2697 21468
rect 2280 21428 2286 21440
rect 2685 21437 2697 21440
rect 2731 21468 2743 21471
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 2731 21440 4905 21468
rect 2731 21437 2743 21440
rect 2685 21431 2743 21437
rect 4893 21437 4905 21440
rect 4939 21437 4951 21471
rect 4893 21431 4951 21437
rect 7190 21428 7196 21480
rect 7248 21428 7254 21480
rect 8297 21471 8355 21477
rect 8297 21437 8309 21471
rect 8343 21437 8355 21471
rect 8297 21431 8355 21437
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 8312 21400 8340 21431
rect 10410 21428 10416 21480
rect 10468 21428 10474 21480
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 10962 21468 10968 21480
rect 10643 21440 10968 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 10962 21428 10968 21440
rect 11020 21428 11026 21480
rect 11974 21428 11980 21480
rect 12032 21468 12038 21480
rect 13173 21471 13231 21477
rect 13173 21468 13185 21471
rect 12032 21440 13185 21468
rect 12032 21428 12038 21440
rect 13173 21437 13185 21440
rect 13219 21437 13231 21471
rect 13173 21431 13231 21437
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21468 13415 21471
rect 13446 21468 13452 21480
rect 13403 21440 13452 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 12066 21400 12072 21412
rect 7616 21372 8340 21400
rect 9600 21372 12072 21400
rect 7616 21360 7622 21372
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 3697 21335 3755 21341
rect 3697 21332 3709 21335
rect 2832 21304 3709 21332
rect 2832 21292 2838 21304
rect 3697 21301 3709 21304
rect 3743 21301 3755 21335
rect 3697 21295 3755 21301
rect 4709 21335 4767 21341
rect 4709 21301 4721 21335
rect 4755 21332 4767 21335
rect 5718 21332 5724 21344
rect 4755 21304 5724 21332
rect 4755 21301 4767 21304
rect 4709 21295 4767 21301
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 9600 21332 9628 21372
rect 12066 21360 12072 21372
rect 12124 21360 12130 21412
rect 14292 21400 14320 21499
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 14976 21508 15669 21536
rect 14976 21496 14982 21508
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 17310 21496 17316 21548
rect 17368 21536 17374 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17368 21508 17509 21536
rect 17368 21496 17374 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 19610 21496 19616 21548
rect 19668 21496 19674 21548
rect 21358 21496 21364 21548
rect 21416 21536 21422 21548
rect 22066 21536 22094 21644
rect 22830 21564 22836 21616
rect 22888 21604 22894 21616
rect 22925 21607 22983 21613
rect 22925 21604 22937 21607
rect 22888 21576 22937 21604
rect 22888 21564 22894 21576
rect 22925 21573 22937 21576
rect 22971 21573 22983 21607
rect 23124 21604 23152 21644
rect 23308 21644 23756 21672
rect 23308 21604 23336 21644
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 23124 21576 23414 21604
rect 22925 21567 22983 21573
rect 21416 21508 22094 21536
rect 21416 21496 21422 21508
rect 22646 21496 22652 21548
rect 22704 21496 22710 21548
rect 14458 21428 14464 21480
rect 14516 21428 14522 21480
rect 22186 21468 22192 21480
rect 20916 21440 22192 21468
rect 19518 21400 19524 21412
rect 14292 21372 19524 21400
rect 19518 21360 19524 21372
rect 19576 21360 19582 21412
rect 6236 21304 9628 21332
rect 6236 21292 6242 21304
rect 9674 21292 9680 21344
rect 9732 21332 9738 21344
rect 9953 21335 10011 21341
rect 9953 21332 9965 21335
rect 9732 21304 9965 21332
rect 9732 21292 9738 21304
rect 9953 21301 9965 21304
rect 9999 21301 10011 21335
rect 9953 21295 10011 21301
rect 12713 21335 12771 21341
rect 12713 21301 12725 21335
rect 12759 21332 12771 21335
rect 13814 21332 13820 21344
rect 12759 21304 13820 21332
rect 12759 21301 12771 21304
rect 12713 21295 12771 21301
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 20916 21332 20944 21440
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 22922 21428 22928 21480
rect 22980 21468 22986 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 22980 21440 24685 21468
rect 22980 21428 22986 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 24673 21431 24731 21437
rect 15519 21304 20944 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 21542 21292 21548 21344
rect 21600 21332 21606 21344
rect 24578 21332 24584 21344
rect 21600 21304 24584 21332
rect 21600 21292 21606 21304
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 2924 21100 3157 21128
rect 2924 21088 2930 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 6546 21088 6552 21140
rect 6604 21128 6610 21140
rect 7653 21131 7711 21137
rect 7653 21128 7665 21131
rect 6604 21100 7665 21128
rect 6604 21088 6610 21100
rect 7653 21097 7665 21100
rect 7699 21097 7711 21131
rect 7653 21091 7711 21097
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 10321 21131 10379 21137
rect 10321 21128 10333 21131
rect 8168 21100 10333 21128
rect 8168 21088 8174 21100
rect 10321 21097 10333 21100
rect 10367 21097 10379 21131
rect 10321 21091 10379 21097
rect 11885 21131 11943 21137
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 11974 21128 11980 21140
rect 11931 21100 11980 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 11974 21088 11980 21100
rect 12032 21088 12038 21140
rect 13722 21088 13728 21140
rect 13780 21088 13786 21140
rect 16666 21128 16672 21140
rect 13832 21100 16672 21128
rect 12618 21060 12624 21072
rect 12544 21032 12624 21060
rect 2774 20952 2780 21004
rect 2832 20952 2838 21004
rect 3970 20952 3976 21004
rect 4028 20952 4034 21004
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 10318 20992 10324 21004
rect 8352 20964 10324 20992
rect 8352 20952 8358 20964
rect 10318 20952 10324 20964
rect 10376 20992 10382 21004
rect 10873 20995 10931 21001
rect 10873 20992 10885 20995
rect 10376 20964 10885 20992
rect 10376 20952 10382 20964
rect 10873 20961 10885 20964
rect 10919 20961 10931 20995
rect 10873 20955 10931 20961
rect 12066 20952 12072 21004
rect 12124 20992 12130 21004
rect 12544 21001 12572 21032
rect 12618 21020 12624 21032
rect 12676 21060 12682 21072
rect 13832 21060 13860 21100
rect 16666 21088 16672 21100
rect 16724 21088 16730 21140
rect 19429 21131 19487 21137
rect 19429 21097 19441 21131
rect 19475 21128 19487 21131
rect 21542 21128 21548 21140
rect 19475 21100 21548 21128
rect 19475 21097 19487 21100
rect 19429 21091 19487 21097
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22370 21088 22376 21140
rect 22428 21088 22434 21140
rect 19334 21060 19340 21072
rect 12676 21032 13860 21060
rect 18800 21032 19340 21060
rect 12676 21020 12682 21032
rect 12345 20995 12403 21001
rect 12345 20992 12357 20995
rect 12124 20964 12357 20992
rect 12124 20952 12130 20964
rect 12345 20961 12357 20964
rect 12391 20961 12403 20995
rect 12345 20955 12403 20961
rect 12529 20995 12587 21001
rect 12529 20961 12541 20995
rect 12575 20961 12587 20995
rect 12529 20955 12587 20961
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 14277 20995 14335 21001
rect 14277 20992 14289 20995
rect 13412 20964 14289 20992
rect 13412 20952 13418 20964
rect 14277 20961 14289 20964
rect 14323 20961 14335 20995
rect 14277 20955 14335 20961
rect 14550 20952 14556 21004
rect 14608 20952 14614 21004
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18800 21001 18828 21032
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 20530 21020 20536 21072
rect 20588 21060 20594 21072
rect 20588 21032 20760 21060
rect 20588 21020 20594 21032
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20961 18843 20995
rect 18785 20955 18843 20961
rect 18966 20952 18972 21004
rect 19024 20992 19030 21004
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 19024 20964 20637 20992
rect 19024 20952 19030 20964
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 20732 20992 20760 21032
rect 23385 20995 23443 21001
rect 23385 20992 23397 20995
rect 20732 20964 23397 20992
rect 20625 20955 20683 20961
rect 23385 20961 23397 20964
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 23474 20952 23480 21004
rect 23532 20952 23538 21004
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2924 20896 2973 20924
rect 2924 20884 2930 20896
rect 2961 20893 2973 20896
rect 3007 20924 3019 20927
rect 3510 20924 3516 20936
rect 3007 20896 3516 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3510 20884 3516 20896
rect 3568 20884 3574 20936
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 11514 20924 11520 20936
rect 10735 20896 11520 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 14182 20924 14188 20936
rect 12299 20896 14188 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 16942 20884 16948 20936
rect 17000 20884 17006 20936
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 17920 20896 18521 20924
rect 17920 20884 17926 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19484 20896 19625 20924
rect 19484 20884 19490 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 22370 20924 22376 20936
rect 22244 20896 22376 20924
rect 22244 20884 22250 20896
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 23293 20927 23351 20933
rect 23293 20924 23305 20927
rect 22796 20896 23305 20924
rect 22796 20884 22802 20896
rect 23293 20893 23305 20896
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 5626 20856 5632 20868
rect 5474 20828 5632 20856
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 7650 20816 7656 20868
rect 7708 20856 7714 20868
rect 8113 20859 8171 20865
rect 8113 20856 8125 20859
rect 7708 20828 8125 20856
rect 7708 20816 7714 20828
rect 8113 20825 8125 20828
rect 8159 20825 8171 20859
rect 16482 20856 16488 20868
rect 15778 20828 16488 20856
rect 8113 20819 8171 20825
rect 16482 20816 16488 20828
rect 16540 20856 16546 20868
rect 17494 20856 17500 20868
rect 16540 20828 17500 20856
rect 16540 20816 16546 20828
rect 17494 20816 17500 20828
rect 17552 20816 17558 20868
rect 20622 20816 20628 20868
rect 20680 20856 20686 20868
rect 20901 20859 20959 20865
rect 20901 20856 20913 20859
rect 20680 20828 20913 20856
rect 20680 20816 20686 20828
rect 20901 20825 20913 20828
rect 20947 20825 20959 20859
rect 21358 20856 21364 20868
rect 20901 20819 20959 20825
rect 21008 20828 21364 20856
rect 5718 20748 5724 20800
rect 5776 20748 5782 20800
rect 6178 20748 6184 20800
rect 6236 20788 6242 20800
rect 6362 20788 6368 20800
rect 6236 20760 6368 20788
rect 6236 20748 6242 20760
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 6454 20748 6460 20800
rect 6512 20788 6518 20800
rect 8021 20791 8079 20797
rect 8021 20788 8033 20791
rect 6512 20760 8033 20788
rect 6512 20748 6518 20760
rect 8021 20757 8033 20760
rect 8067 20788 8079 20791
rect 8570 20788 8576 20800
rect 8067 20760 8576 20788
rect 8067 20757 8079 20760
rect 8021 20751 8079 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9214 20748 9220 20800
rect 9272 20788 9278 20800
rect 10686 20788 10692 20800
rect 9272 20760 10692 20788
rect 9272 20748 9278 20760
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 10781 20791 10839 20797
rect 10781 20757 10793 20791
rect 10827 20788 10839 20791
rect 11606 20788 11612 20800
rect 10827 20760 11612 20788
rect 10827 20757 10839 20760
rect 10781 20751 10839 20757
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 16022 20748 16028 20800
rect 16080 20748 16086 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 16632 20760 18153 20788
rect 16632 20748 16638 20760
rect 18141 20757 18153 20760
rect 18187 20757 18199 20791
rect 18141 20751 18199 20757
rect 20346 20748 20352 20800
rect 20404 20788 20410 20800
rect 21008 20788 21036 20828
rect 21358 20816 21364 20828
rect 21416 20816 21422 20868
rect 20404 20760 21036 20788
rect 20404 20748 20410 20760
rect 22922 20748 22928 20800
rect 22980 20748 22986 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 7377 20587 7435 20593
rect 7377 20553 7389 20587
rect 7423 20584 7435 20587
rect 7742 20584 7748 20596
rect 7423 20556 7748 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 12069 20587 12127 20593
rect 12069 20553 12081 20587
rect 12115 20584 12127 20587
rect 12158 20584 12164 20596
rect 12115 20556 12164 20584
rect 12115 20553 12127 20556
rect 12069 20547 12127 20553
rect 12158 20544 12164 20556
rect 12216 20544 12222 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14737 20587 14795 20593
rect 14737 20584 14749 20587
rect 13872 20556 14749 20584
rect 13872 20544 13878 20556
rect 14737 20553 14749 20556
rect 14783 20553 14795 20587
rect 14737 20547 14795 20553
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 15102 20584 15108 20596
rect 14875 20556 15108 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17221 20587 17279 20593
rect 17221 20584 17233 20587
rect 17000 20556 17233 20584
rect 17000 20544 17006 20556
rect 17221 20553 17233 20556
rect 17267 20553 17279 20587
rect 17221 20547 17279 20553
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20584 17371 20587
rect 17402 20584 17408 20596
rect 17359 20556 17408 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 22373 20587 22431 20593
rect 22373 20553 22385 20587
rect 22419 20584 22431 20587
rect 22922 20584 22928 20596
rect 22419 20556 22928 20584
rect 22419 20553 22431 20556
rect 22373 20547 22431 20553
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 23474 20544 23480 20596
rect 23532 20584 23538 20596
rect 23532 20556 23704 20584
rect 23532 20544 23538 20556
rect 6822 20476 6828 20528
rect 6880 20516 6886 20528
rect 18966 20516 18972 20528
rect 6880 20488 9338 20516
rect 18800 20488 18972 20516
rect 6880 20476 6886 20488
rect 1762 20408 1768 20460
rect 1820 20408 1826 20460
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7742 20448 7748 20460
rect 7156 20420 7748 20448
rect 7156 20408 7162 20420
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 8573 20451 8631 20457
rect 8573 20448 8585 20451
rect 8076 20420 8585 20448
rect 8076 20408 8082 20420
rect 8573 20417 8585 20420
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 17034 20448 17040 20460
rect 15795 20420 17040 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 18800 20457 18828 20488
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 20346 20516 20352 20528
rect 20286 20488 20352 20516
rect 20346 20476 20352 20488
rect 20404 20476 20410 20528
rect 20806 20476 20812 20528
rect 20864 20516 20870 20528
rect 21269 20519 21327 20525
rect 21269 20516 21281 20519
rect 20864 20488 21281 20516
rect 20864 20476 20870 20488
rect 21269 20485 21281 20488
rect 21315 20485 21327 20519
rect 21269 20479 21327 20485
rect 22465 20519 22523 20525
rect 22465 20485 22477 20519
rect 22511 20516 22523 20519
rect 22554 20516 22560 20528
rect 22511 20488 22560 20516
rect 22511 20485 22523 20488
rect 22465 20479 22523 20485
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 23676 20525 23704 20556
rect 23661 20519 23719 20525
rect 23661 20485 23673 20519
rect 23707 20485 23719 20519
rect 23661 20479 23719 20485
rect 23750 20476 23756 20528
rect 23808 20516 23814 20528
rect 23808 20488 24150 20516
rect 23808 20476 23814 20488
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 23385 20451 23443 20457
rect 23385 20448 23397 20451
rect 22704 20420 23397 20448
rect 22704 20408 22710 20420
rect 23385 20417 23397 20420
rect 23431 20417 23443 20451
rect 23385 20411 23443 20417
rect 1302 20340 1308 20392
rect 1360 20380 1366 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1360 20352 2053 20380
rect 1360 20340 1366 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 7852 20312 7880 20343
rect 7926 20340 7932 20392
rect 7984 20340 7990 20392
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20380 8907 20383
rect 12066 20380 12072 20392
rect 8895 20352 12072 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 12158 20340 12164 20392
rect 12216 20340 12222 20392
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 8570 20312 8576 20324
rect 7852 20284 8576 20312
rect 8570 20272 8576 20284
rect 8628 20272 8634 20324
rect 10134 20272 10140 20324
rect 10192 20312 10198 20324
rect 11054 20312 11060 20324
rect 10192 20284 11060 20312
rect 10192 20272 10198 20284
rect 11054 20272 11060 20284
rect 11112 20312 11118 20324
rect 12268 20312 12296 20343
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14458 20380 14464 20392
rect 13504 20352 14464 20380
rect 13504 20340 13510 20352
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 16022 20380 16028 20392
rect 15059 20352 16028 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20380 17555 20383
rect 18506 20380 18512 20392
rect 17543 20352 18512 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 18506 20340 18512 20352
rect 18564 20380 18570 20392
rect 19061 20383 19119 20389
rect 19061 20380 19073 20383
rect 18564 20352 19073 20380
rect 18564 20340 18570 20352
rect 19061 20349 19073 20352
rect 19107 20349 19119 20383
rect 19061 20343 19119 20349
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 11112 20284 12296 20312
rect 11112 20272 11118 20284
rect 20622 20272 20628 20324
rect 20680 20312 20686 20324
rect 21453 20315 21511 20321
rect 20680 20284 20852 20312
rect 20680 20272 20686 20284
rect 11146 20204 11152 20256
rect 11204 20204 11210 20256
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 11701 20247 11759 20253
rect 11701 20244 11713 20247
rect 11296 20216 11713 20244
rect 11296 20204 11302 20216
rect 11701 20213 11713 20216
rect 11747 20213 11759 20247
rect 11701 20207 11759 20213
rect 14369 20247 14427 20253
rect 14369 20213 14381 20247
rect 14415 20244 14427 20247
rect 14734 20244 14740 20256
rect 14415 20216 14740 20244
rect 14415 20213 14427 20216
rect 14369 20207 14427 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 15565 20247 15623 20253
rect 15565 20213 15577 20247
rect 15611 20244 15623 20247
rect 15838 20244 15844 20256
rect 15611 20216 15844 20244
rect 15611 20213 15623 20216
rect 15565 20207 15623 20213
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 16853 20247 16911 20253
rect 16853 20213 16865 20247
rect 16899 20244 16911 20247
rect 18230 20244 18236 20256
rect 16899 20216 18236 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 20533 20247 20591 20253
rect 20533 20213 20545 20247
rect 20579 20244 20591 20247
rect 20714 20244 20720 20256
rect 20579 20216 20720 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 20824 20244 20852 20284
rect 21453 20281 21465 20315
rect 21499 20312 21511 20315
rect 21634 20312 21640 20324
rect 21499 20284 21640 20312
rect 21499 20281 21511 20284
rect 21453 20275 21511 20281
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 20824 20216 22017 20244
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22572 20244 22600 20343
rect 22830 20244 22836 20256
rect 22572 20216 22836 20244
rect 22005 20207 22063 20213
rect 22830 20204 22836 20216
rect 22888 20244 22894 20256
rect 25133 20247 25191 20253
rect 25133 20244 25145 20247
rect 22888 20216 25145 20244
rect 22888 20204 22894 20216
rect 25133 20213 25145 20216
rect 25179 20213 25191 20247
rect 25133 20207 25191 20213
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 7006 20040 7012 20052
rect 6012 20012 7012 20040
rect 4617 19907 4675 19913
rect 4617 19873 4629 19907
rect 4663 19904 4675 19907
rect 6012 19904 6040 20012
rect 7006 20000 7012 20012
rect 7064 20040 7070 20052
rect 7064 20012 7880 20040
rect 7064 20000 7070 20012
rect 4663 19876 6040 19904
rect 6089 19907 6147 19913
rect 4663 19873 4675 19876
rect 4617 19867 4675 19873
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6825 19907 6883 19913
rect 6825 19904 6837 19907
rect 6135 19876 6837 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6825 19873 6837 19876
rect 6871 19904 6883 19907
rect 7190 19904 7196 19916
rect 6871 19876 7196 19904
rect 6871 19873 6883 19876
rect 6825 19867 6883 19873
rect 7190 19864 7196 19876
rect 7248 19864 7254 19916
rect 7852 19904 7880 20012
rect 9122 20000 9128 20052
rect 9180 20000 9186 20052
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 12894 20040 12900 20052
rect 12400 20012 12900 20040
rect 12400 20000 12406 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 21910 20040 21916 20052
rect 16071 20012 21916 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 20714 19972 20720 19984
rect 18616 19944 20720 19972
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 7852 19876 9689 19904
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 11238 19904 11244 19916
rect 9677 19867 9735 19873
rect 10612 19876 11244 19904
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 3326 19836 3332 19848
rect 2271 19808 3332 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19805 4399 19839
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 4341 19799 4399 19805
rect 6012 19808 6561 19836
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 2041 19703 2099 19709
rect 2041 19700 2053 19703
rect 1912 19672 2053 19700
rect 1912 19660 1918 19672
rect 2041 19669 2053 19672
rect 2087 19669 2099 19703
rect 4356 19700 4384 19799
rect 5626 19728 5632 19780
rect 5684 19728 5690 19780
rect 5442 19700 5448 19712
rect 4356 19672 5448 19700
rect 2041 19663 2099 19669
rect 5442 19660 5448 19672
rect 5500 19700 5506 19712
rect 6012 19700 6040 19808
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 10612 19836 10640 19876
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 11793 19907 11851 19913
rect 11793 19904 11805 19907
rect 11388 19876 11805 19904
rect 11388 19864 11394 19876
rect 11793 19873 11805 19876
rect 11839 19873 11851 19907
rect 11793 19867 11851 19873
rect 9539 19808 10640 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 11146 19796 11152 19848
rect 11204 19836 11210 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11204 19808 11713 19836
rect 11204 19796 11210 19808
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 11808 19836 11836 19867
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 18414 19864 18420 19916
rect 18472 19864 18478 19916
rect 18616 19913 18644 19944
rect 20714 19932 20720 19944
rect 20772 19932 20778 19984
rect 22646 19972 22652 19984
rect 21560 19944 22652 19972
rect 21560 19913 21588 19944
rect 22646 19932 22652 19944
rect 22704 19932 22710 19984
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 13354 19836 13360 19848
rect 11808 19808 13360 19836
rect 11701 19799 11759 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 14918 19796 14924 19848
rect 14976 19836 14982 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 14976 19808 16221 19836
rect 14976 19796 14982 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 17310 19796 17316 19848
rect 17368 19796 17374 19848
rect 18322 19796 18328 19848
rect 18380 19836 18386 19848
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 18380 19808 20729 19836
rect 18380 19796 18386 19808
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 25222 19836 25228 19848
rect 22879 19808 25228 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 25222 19796 25228 19808
rect 25280 19796 25286 19848
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 6822 19768 6828 19780
rect 6236 19740 6828 19768
rect 6236 19728 6242 19740
rect 6822 19728 6828 19740
rect 6880 19768 6886 19780
rect 8573 19771 8631 19777
rect 6880 19740 7314 19768
rect 6880 19728 6886 19740
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 8619 19740 11744 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 11716 19712 11744 19740
rect 17494 19728 17500 19780
rect 17552 19728 17558 19780
rect 18598 19768 18604 19780
rect 17972 19740 18604 19768
rect 5500 19672 6040 19700
rect 9585 19703 9643 19709
rect 5500 19660 5506 19672
rect 9585 19669 9597 19703
rect 9631 19700 9643 19703
rect 10134 19700 10140 19712
rect 9631 19672 10140 19700
rect 9631 19669 9643 19672
rect 9585 19663 9643 19669
rect 10134 19660 10140 19672
rect 10192 19660 10198 19712
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 11333 19703 11391 19709
rect 11333 19700 11345 19703
rect 11204 19672 11345 19700
rect 11204 19660 11210 19672
rect 11333 19669 11345 19672
rect 11379 19669 11391 19703
rect 11333 19663 11391 19669
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 12250 19700 12256 19712
rect 11756 19672 12256 19700
rect 11756 19660 11762 19672
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 17972 19709 18000 19740
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 20073 19771 20131 19777
rect 20073 19768 20085 19771
rect 19300 19740 20085 19768
rect 19300 19728 19306 19740
rect 20073 19737 20085 19740
rect 20119 19737 20131 19771
rect 20073 19731 20131 19737
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 21818 19768 21824 19780
rect 20303 19740 21824 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19669 18015 19703
rect 17957 19663 18015 19669
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18325 19703 18383 19709
rect 18325 19700 18337 19703
rect 18288 19672 18337 19700
rect 18288 19660 18294 19672
rect 18325 19669 18337 19672
rect 18371 19669 18383 19703
rect 18325 19663 18383 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 4798 19456 4804 19508
rect 4856 19456 4862 19508
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7524 19468 8125 19496
rect 7524 19456 7530 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 8573 19499 8631 19505
rect 8573 19465 8585 19499
rect 8619 19496 8631 19499
rect 9674 19496 9680 19508
rect 8619 19468 9680 19496
rect 8619 19465 8631 19468
rect 8573 19459 8631 19465
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 10284 19468 10425 19496
rect 10284 19456 10290 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 11054 19496 11060 19508
rect 10413 19459 10471 19465
rect 10796 19468 11060 19496
rect 7834 19388 7840 19440
rect 7892 19428 7898 19440
rect 10796 19428 10824 19468
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 11664 19468 13093 19496
rect 11664 19456 11670 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 13081 19459 13139 19465
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 17865 19499 17923 19505
rect 15988 19468 17356 19496
rect 15988 19456 15994 19468
rect 7892 19400 10824 19428
rect 10873 19431 10931 19437
rect 7892 19388 7898 19400
rect 10873 19397 10885 19431
rect 10919 19428 10931 19431
rect 11790 19428 11796 19440
rect 10919 19400 11796 19428
rect 10919 19397 10931 19400
rect 10873 19391 10931 19397
rect 11790 19388 11796 19400
rect 11848 19388 11854 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 13449 19431 13507 19437
rect 12124 19400 12480 19428
rect 12124 19388 12130 19400
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19360 5043 19363
rect 7558 19360 7564 19372
rect 5031 19332 7564 19360
rect 5031 19329 5043 19332
rect 4985 19323 5043 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8478 19320 8484 19372
rect 8536 19320 8542 19372
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19360 10839 19363
rect 11698 19360 11704 19372
rect 10827 19332 11704 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19292 8815 19295
rect 9398 19292 9404 19304
rect 8803 19264 9404 19292
rect 8803 19261 8815 19264
rect 8757 19255 8815 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10376 19264 10977 19292
rect 10376 19252 10382 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 12452 19292 12480 19400
rect 13449 19397 13461 19431
rect 13495 19428 13507 19431
rect 17034 19428 17040 19440
rect 13495 19400 17040 19428
rect 13495 19397 13507 19400
rect 13449 19391 13507 19397
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 17218 19388 17224 19440
rect 17276 19388 17282 19440
rect 17328 19428 17356 19468
rect 17865 19465 17877 19499
rect 17911 19496 17923 19499
rect 20990 19496 20996 19508
rect 17911 19468 20996 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 19429 19431 19487 19437
rect 19429 19428 19441 19431
rect 17328 19400 19441 19428
rect 19429 19397 19441 19400
rect 19475 19397 19487 19431
rect 19429 19391 19487 19397
rect 21269 19431 21327 19437
rect 21269 19397 21281 19431
rect 21315 19428 21327 19431
rect 22186 19428 22192 19440
rect 21315 19400 22192 19428
rect 21315 19397 21327 19400
rect 21269 19391 21327 19397
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23293 19431 23351 19437
rect 23293 19397 23305 19431
rect 23339 19428 23351 19431
rect 24854 19428 24860 19440
rect 23339 19400 24860 19428
rect 23339 19397 23351 19400
rect 23293 19391 23351 19397
rect 24854 19388 24860 19400
rect 24912 19388 24918 19440
rect 13538 19320 13544 19372
rect 13596 19320 13602 19372
rect 15286 19320 15292 19372
rect 15344 19360 15350 19372
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 15344 19332 18061 19360
rect 15344 19320 15350 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 21082 19360 21088 19372
rect 20303 19332 21088 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 22094 19320 22100 19372
rect 22152 19320 22158 19372
rect 24121 19363 24179 19369
rect 24121 19329 24133 19363
rect 24167 19360 24179 19363
rect 25038 19360 25044 19372
rect 24167 19332 25044 19360
rect 24167 19329 24179 19332
rect 24121 19323 24179 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 12618 19292 12624 19304
rect 12452 19264 12624 19292
rect 10965 19255 11023 19261
rect 12618 19252 12624 19264
rect 12676 19292 12682 19304
rect 13633 19295 13691 19301
rect 13633 19292 13645 19295
rect 12676 19264 13645 19292
rect 12676 19252 12682 19264
rect 13633 19261 13645 19264
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 24670 19252 24676 19304
rect 24728 19252 24734 19304
rect 19613 19227 19671 19233
rect 19613 19193 19625 19227
rect 19659 19224 19671 19227
rect 23474 19224 23480 19236
rect 19659 19196 23480 19224
rect 19659 19193 19671 19196
rect 19613 19187 19671 19193
rect 23474 19184 23480 19196
rect 23532 19184 23538 19236
rect 5626 19116 5632 19168
rect 5684 19156 5690 19168
rect 6178 19156 6184 19168
rect 5684 19128 6184 19156
rect 5684 19116 5690 19128
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 12894 19156 12900 19168
rect 11388 19128 12900 19156
rect 11388 19116 11394 19128
rect 12894 19116 12900 19128
rect 12952 19156 12958 19168
rect 14458 19156 14464 19168
rect 12952 19128 14464 19156
rect 12952 19116 12958 19128
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 17092 19128 17325 19156
rect 17092 19116 17098 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18966 19156 18972 19168
rect 18555 19128 18972 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 20438 19156 20444 19168
rect 20312 19128 20444 19156
rect 20312 19116 20318 19128
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22370 19156 22376 19168
rect 22152 19128 22376 19156
rect 22152 19116 22158 19128
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 3786 18912 3792 18964
rect 3844 18952 3850 18964
rect 3973 18955 4031 18961
rect 3973 18952 3985 18955
rect 3844 18924 3985 18952
rect 3844 18912 3850 18924
rect 3973 18921 3985 18924
rect 4019 18921 4031 18955
rect 3973 18915 4031 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7064 18924 7205 18952
rect 7064 18912 7070 18924
rect 7193 18921 7205 18924
rect 7239 18921 7251 18955
rect 7193 18915 7251 18921
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 8628 18924 10701 18952
rect 8628 18912 8634 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 11020 18924 13400 18952
rect 11020 18912 11026 18924
rect 3418 18776 3424 18828
rect 3476 18816 3482 18828
rect 7742 18816 7748 18828
rect 3476 18788 7748 18816
rect 3476 18776 3482 18788
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 11330 18776 11336 18828
rect 11388 18776 11394 18828
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 12802 18816 12808 18828
rect 11664 18788 12808 18816
rect 11664 18776 11670 18788
rect 12802 18776 12808 18788
rect 12860 18816 12866 18828
rect 13372 18825 13400 18924
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 20438 18884 20444 18896
rect 17267 18856 20444 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 20438 18844 20444 18856
rect 20496 18844 20502 18896
rect 20993 18887 21051 18893
rect 20993 18853 21005 18887
rect 21039 18884 21051 18887
rect 22186 18884 22192 18896
rect 21039 18856 22192 18884
rect 21039 18853 21051 18856
rect 20993 18847 21051 18853
rect 22186 18844 22192 18856
rect 22244 18844 22250 18896
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 12860 18788 13185 18816
rect 12860 18776 12866 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13173 18779 13231 18785
rect 13357 18819 13415 18825
rect 13357 18785 13369 18819
rect 13403 18816 13415 18819
rect 13446 18816 13452 18828
rect 13403 18788 13452 18816
rect 13403 18785 13415 18788
rect 13357 18779 13415 18785
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17184 18788 17693 18816
rect 17184 18776 17190 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18816 17923 18819
rect 19242 18816 19248 18828
rect 17911 18788 19248 18816
rect 17911 18785 17923 18788
rect 17865 18779 17923 18785
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19886 18776 19892 18828
rect 19944 18776 19950 18828
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18816 20131 18819
rect 21358 18816 21364 18828
rect 20119 18788 21364 18816
rect 20119 18785 20131 18788
rect 20073 18779 20131 18785
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 22554 18816 22560 18828
rect 21683 18788 22560 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 22554 18776 22560 18788
rect 22612 18816 22618 18828
rect 23937 18819 23995 18825
rect 23937 18816 23949 18819
rect 22612 18788 23949 18816
rect 22612 18776 22618 18788
rect 23937 18785 23949 18788
rect 23983 18785 23995 18819
rect 23937 18779 23995 18785
rect 2222 18708 2228 18760
rect 2280 18708 2286 18760
rect 4154 18708 4160 18760
rect 4212 18708 4218 18760
rect 5442 18708 5448 18760
rect 5500 18708 5506 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 12710 18748 12716 18760
rect 11103 18720 12716 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 12710 18708 12716 18720
rect 12768 18748 12774 18760
rect 14182 18748 14188 18760
rect 12768 18720 14188 18748
rect 12768 18708 12774 18720
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 16574 18708 16580 18760
rect 16632 18708 16638 18760
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 19797 18751 19855 18757
rect 19797 18748 19809 18751
rect 18564 18720 19809 18748
rect 18564 18708 18570 18720
rect 19797 18717 19809 18720
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 21726 18748 21732 18760
rect 21499 18720 21732 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22060 18720 22201 18748
rect 22060 18708 22066 18720
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 24673 18751 24731 18757
rect 24673 18748 24685 18751
rect 24636 18720 24685 18748
rect 24636 18708 24642 18720
rect 24673 18717 24685 18720
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 5721 18683 5779 18689
rect 5721 18649 5733 18683
rect 5767 18649 5779 18683
rect 5721 18643 5779 18649
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 2041 18615 2099 18621
rect 2041 18612 2053 18615
rect 1820 18584 2053 18612
rect 1820 18572 1826 18584
rect 2041 18581 2053 18584
rect 2087 18581 2099 18615
rect 5736 18612 5764 18643
rect 6178 18640 6184 18692
rect 6236 18640 6242 18692
rect 12342 18680 12348 18692
rect 11256 18652 12348 18680
rect 11256 18624 11284 18652
rect 12342 18640 12348 18652
rect 12400 18640 12406 18692
rect 13538 18640 13544 18692
rect 13596 18680 13602 18692
rect 17589 18683 17647 18689
rect 17589 18680 17601 18683
rect 13596 18652 17601 18680
rect 13596 18640 13602 18652
rect 17589 18649 17601 18652
rect 17635 18649 17647 18683
rect 17589 18643 17647 18649
rect 19058 18640 19064 18692
rect 19116 18680 19122 18692
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 19116 18652 21373 18680
rect 19116 18640 19122 18652
rect 21361 18649 21373 18652
rect 21407 18649 21419 18683
rect 21361 18643 21419 18649
rect 22465 18683 22523 18689
rect 22465 18649 22477 18683
rect 22511 18649 22523 18683
rect 23750 18680 23756 18692
rect 23690 18652 23756 18680
rect 22465 18643 22523 18649
rect 7834 18612 7840 18624
rect 5736 18584 7840 18612
rect 2041 18575 2099 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 11149 18615 11207 18621
rect 11149 18581 11161 18615
rect 11195 18612 11207 18615
rect 11238 18612 11244 18624
rect 11195 18584 11244 18612
rect 11195 18581 11207 18584
rect 11149 18575 11207 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12713 18615 12771 18621
rect 12713 18612 12725 18615
rect 12124 18584 12725 18612
rect 12124 18572 12130 18584
rect 12713 18581 12725 18584
rect 12759 18581 12771 18615
rect 12713 18575 12771 18581
rect 13081 18615 13139 18621
rect 13081 18581 13093 18615
rect 13127 18612 13139 18615
rect 15930 18612 15936 18624
rect 13127 18584 15936 18612
rect 13127 18581 13139 18584
rect 13081 18575 13139 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 16669 18615 16727 18621
rect 16669 18612 16681 18615
rect 16632 18584 16681 18612
rect 16632 18572 16638 18584
rect 16669 18581 16681 18584
rect 16715 18581 16727 18615
rect 16669 18575 16727 18581
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 20162 18612 20168 18624
rect 19475 18584 20168 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 22480 18612 22508 18643
rect 23750 18640 23756 18652
rect 23808 18640 23814 18692
rect 22646 18612 22652 18624
rect 22480 18584 22652 18612
rect 22646 18572 22652 18584
rect 22704 18612 22710 18624
rect 23290 18612 23296 18624
rect 22704 18584 23296 18612
rect 22704 18572 22710 18584
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 24210 18572 24216 18624
rect 24268 18612 24274 18624
rect 24765 18615 24823 18621
rect 24765 18612 24777 18615
rect 24268 18584 24777 18612
rect 24268 18572 24274 18584
rect 24765 18581 24777 18584
rect 24811 18581 24823 18615
rect 24765 18575 24823 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 10594 18408 10600 18420
rect 9232 18380 10600 18408
rect 6178 18300 6184 18352
rect 6236 18340 6242 18352
rect 6236 18312 7682 18340
rect 6236 18300 6242 18312
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 1854 18272 1860 18284
rect 1811 18244 1860 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1360 18176 2053 18204
rect 1360 18164 1366 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 6914 18164 6920 18216
rect 6972 18164 6978 18216
rect 7193 18207 7251 18213
rect 7193 18173 7205 18207
rect 7239 18204 7251 18207
rect 9232 18204 9260 18380
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 11054 18368 11060 18420
rect 11112 18368 11118 18420
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 11756 18380 12449 18408
rect 11756 18368 11762 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 12805 18411 12863 18417
rect 12805 18377 12817 18411
rect 12851 18408 12863 18411
rect 13538 18408 13544 18420
rect 12851 18380 13544 18408
rect 12851 18377 12863 18380
rect 12805 18371 12863 18377
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 20898 18408 20904 18420
rect 19628 18380 20904 18408
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 9732 18312 10074 18340
rect 9732 18300 9738 18312
rect 10870 18300 10876 18352
rect 10928 18340 10934 18352
rect 12342 18340 12348 18352
rect 10928 18312 12348 18340
rect 10928 18300 10934 18312
rect 12342 18300 12348 18312
rect 12400 18340 12406 18352
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 12400 18312 14105 18340
rect 12400 18300 12406 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 14093 18303 14151 18309
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18340 18107 18343
rect 18322 18340 18328 18352
rect 18095 18312 18328 18340
rect 18095 18309 18107 18312
rect 18049 18303 18107 18309
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 13722 18272 13728 18284
rect 12943 18244 13728 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 18966 18272 18972 18284
rect 14047 18244 18972 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 19628 18281 19656 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 23290 18368 23296 18420
rect 23348 18408 23354 18420
rect 24489 18411 24547 18417
rect 24489 18408 24501 18411
rect 23348 18380 24501 18408
rect 23348 18368 23354 18380
rect 24489 18377 24501 18380
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 22462 18340 22468 18352
rect 20272 18312 22468 18340
rect 20272 18281 20300 18312
rect 22462 18300 22468 18312
rect 22520 18300 22526 18352
rect 22738 18300 22744 18352
rect 22796 18340 22802 18352
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 22796 18312 23029 18340
rect 22796 18300 22802 18312
rect 23017 18309 23029 18312
rect 23063 18309 23075 18343
rect 23017 18303 23075 18309
rect 23750 18300 23756 18352
rect 23808 18300 23814 18352
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 22370 18272 22376 18284
rect 22244 18244 22376 18272
rect 22244 18232 22250 18244
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 7239 18176 9260 18204
rect 9309 18207 9367 18213
rect 7239 18173 7251 18176
rect 7193 18167 7251 18173
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 11330 18204 11336 18216
rect 9631 18176 11336 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8665 18071 8723 18077
rect 8665 18068 8677 18071
rect 7892 18040 8677 18068
rect 7892 18028 7898 18040
rect 8665 18037 8677 18040
rect 8711 18037 8723 18071
rect 9324 18068 9352 18167
rect 11330 18164 11336 18176
rect 11388 18164 11394 18216
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12989 18207 13047 18213
rect 12989 18204 13001 18207
rect 12676 18176 13001 18204
rect 12676 18164 12682 18176
rect 12989 18173 13001 18176
rect 13035 18173 13047 18207
rect 12989 18167 13047 18173
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14458 18204 14464 18216
rect 14323 18176 14464 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 17460 18176 18797 18204
rect 17460 18164 17466 18176
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 21269 18207 21327 18213
rect 21269 18173 21281 18207
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 12158 18096 12164 18148
rect 12216 18136 12222 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 12216 18108 13645 18136
rect 12216 18096 12222 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 21284 18136 21312 18167
rect 22002 18164 22008 18216
rect 22060 18204 22066 18216
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22060 18176 22753 18204
rect 22060 18164 22066 18176
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 22741 18167 22799 18173
rect 21284 18108 22324 18136
rect 13633 18099 13691 18105
rect 10226 18068 10232 18080
rect 9324 18040 10232 18068
rect 8665 18031 8723 18037
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 16574 18068 16580 18080
rect 13596 18040 16580 18068
rect 13596 18028 13602 18040
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 20070 18068 20076 18080
rect 19475 18040 20076 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 22186 18028 22192 18080
rect 22244 18028 22250 18080
rect 22296 18068 22324 18108
rect 22462 18096 22468 18148
rect 22520 18136 22526 18148
rect 22646 18136 22652 18148
rect 22520 18108 22652 18136
rect 22520 18096 22526 18108
rect 22646 18096 22652 18108
rect 22704 18096 22710 18148
rect 23382 18068 23388 18080
rect 22296 18040 23388 18068
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 4430 17824 4436 17876
rect 4488 17864 4494 17876
rect 9401 17867 9459 17873
rect 4488 17836 9168 17864
rect 4488 17824 4494 17836
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 5442 17728 5448 17740
rect 4847 17700 5448 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 6178 17620 6184 17672
rect 6236 17620 6242 17672
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 9140 17669 9168 17836
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 11514 17864 11520 17876
rect 9447 17836 11520 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 17681 17867 17739 17873
rect 17681 17864 17693 17867
rect 16724 17836 17693 17864
rect 16724 17824 16730 17836
rect 17681 17833 17693 17836
rect 17727 17833 17739 17867
rect 17681 17827 17739 17833
rect 18782 17824 18788 17876
rect 18840 17864 18846 17876
rect 19334 17864 19340 17876
rect 18840 17836 19340 17864
rect 18840 17824 18846 17836
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20254 17864 20260 17876
rect 19444 17836 20260 17864
rect 18414 17756 18420 17808
rect 18472 17796 18478 17808
rect 19444 17796 19472 17836
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 18472 17768 19472 17796
rect 18472 17756 18478 17768
rect 18800 17740 18828 17768
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12032 17700 13093 17728
rect 12032 17688 12038 17700
rect 13081 17697 13093 17700
rect 13127 17728 13139 17731
rect 13538 17728 13544 17740
rect 13127 17700 13544 17728
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15470 17728 15476 17740
rect 14967 17700 15476 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15933 17731 15991 17737
rect 15933 17697 15945 17731
rect 15979 17728 15991 17731
rect 17402 17728 17408 17740
rect 15979 17700 17408 17728
rect 15979 17697 15991 17700
rect 15933 17691 15991 17697
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 18782 17688 18788 17740
rect 18840 17688 18846 17740
rect 19242 17688 19248 17740
rect 19300 17728 19306 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19300 17700 19717 17728
rect 19300 17688 19306 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 20404 17700 20760 17728
rect 20404 17688 20410 17700
rect 8389 17663 8447 17669
rect 8389 17660 8401 17663
rect 6972 17632 8401 17660
rect 6972 17620 6978 17632
rect 8389 17629 8401 17632
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17660 13047 17663
rect 14274 17660 14280 17672
rect 13035 17632 14280 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 17310 17620 17316 17672
rect 17368 17620 17374 17672
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 19150 17660 19156 17672
rect 18371 17632 19156 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 20732 17604 20760 17700
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 22278 17620 22284 17672
rect 22336 17660 22342 17672
rect 22649 17663 22707 17669
rect 22649 17660 22661 17663
rect 22336 17632 22661 17660
rect 22336 17620 22342 17632
rect 22649 17629 22661 17632
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17561 5135 17595
rect 7282 17592 7288 17604
rect 5077 17555 5135 17561
rect 6472 17564 7288 17592
rect 5092 17524 5120 17555
rect 6472 17524 6500 17564
rect 7282 17552 7288 17564
rect 7340 17552 7346 17604
rect 7653 17595 7711 17601
rect 7653 17561 7665 17595
rect 7699 17592 7711 17595
rect 10042 17592 10048 17604
rect 7699 17564 10048 17592
rect 7699 17561 7711 17564
rect 7653 17555 7711 17561
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 10226 17552 10232 17604
rect 10284 17592 10290 17604
rect 10781 17595 10839 17601
rect 10781 17592 10793 17595
rect 10284 17564 10793 17592
rect 10284 17552 10290 17564
rect 10781 17561 10793 17564
rect 10827 17561 10839 17595
rect 10781 17555 10839 17561
rect 12897 17595 12955 17601
rect 12897 17561 12909 17595
rect 12943 17592 12955 17595
rect 16209 17595 16267 17601
rect 12943 17564 14320 17592
rect 12943 17561 12955 17564
rect 12897 17555 12955 17561
rect 5092 17496 6500 17524
rect 6546 17484 6552 17536
rect 6604 17484 6610 17536
rect 9582 17484 9588 17536
rect 9640 17484 9646 17536
rect 12526 17484 12532 17536
rect 12584 17484 12590 17536
rect 14292 17533 14320 17564
rect 16209 17561 16221 17595
rect 16255 17561 16267 17595
rect 18690 17592 18696 17604
rect 16209 17555 16267 17561
rect 17604 17564 18696 17592
rect 14277 17527 14335 17533
rect 14277 17493 14289 17527
rect 14323 17493 14335 17527
rect 14277 17487 14335 17493
rect 14642 17484 14648 17536
rect 14700 17484 14706 17536
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 15102 17524 15108 17536
rect 14783 17496 15108 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 16224 17524 16252 17555
rect 17604 17524 17632 17564
rect 18690 17552 18696 17564
rect 18748 17552 18754 17604
rect 20714 17552 20720 17604
rect 20772 17552 20778 17604
rect 16224 17496 17632 17524
rect 18417 17527 18475 17533
rect 18417 17493 18429 17527
rect 18463 17524 18475 17527
rect 19702 17524 19708 17536
rect 18463 17496 19708 17524
rect 18463 17493 18475 17496
rect 18417 17487 18475 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 20530 17524 20536 17536
rect 20036 17496 20536 17524
rect 20036 17484 20042 17496
rect 20530 17484 20536 17496
rect 20588 17524 20594 17536
rect 21177 17527 21235 17533
rect 21177 17524 21189 17527
rect 20588 17496 21189 17524
rect 20588 17484 20594 17496
rect 21177 17493 21189 17496
rect 21223 17493 21235 17527
rect 21177 17487 21235 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 4212 17292 5273 17320
rect 4212 17280 4218 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 5721 17323 5779 17329
rect 5721 17289 5733 17323
rect 5767 17320 5779 17323
rect 8665 17323 8723 17329
rect 8665 17320 8677 17323
rect 5767 17292 8677 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 8665 17289 8677 17292
rect 8711 17289 8723 17323
rect 8665 17283 8723 17289
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9171 17292 10088 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 5166 17212 5172 17264
rect 5224 17252 5230 17264
rect 5224 17224 7144 17252
rect 5224 17212 5230 17224
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 7006 17184 7012 17196
rect 5675 17156 7012 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 7116 17184 7144 17224
rect 7282 17212 7288 17264
rect 7340 17252 7346 17264
rect 9033 17255 9091 17261
rect 7340 17224 8984 17252
rect 7340 17212 7346 17224
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7116 17156 7849 17184
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8956 17184 8984 17224
rect 9033 17221 9045 17255
rect 9079 17252 9091 17255
rect 9079 17224 9996 17252
rect 9079 17221 9091 17224
rect 9033 17215 9091 17221
rect 7975 17156 8892 17184
rect 8956 17156 9260 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6546 17116 6552 17128
rect 5951 17088 6552 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8036 17048 8064 17079
rect 7892 17020 8064 17048
rect 8864 17048 8892 17156
rect 9232 17125 9260 17156
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17085 9275 17119
rect 9217 17079 9275 17085
rect 9858 17048 9864 17060
rect 8864 17020 9864 17048
rect 7892 17008 7898 17020
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 7469 16983 7527 16989
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 9306 16980 9312 16992
rect 7515 16952 9312 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9968 16980 9996 17224
rect 10060 17184 10088 17292
rect 10134 17280 10140 17332
rect 10192 17280 10198 17332
rect 12066 17280 12072 17332
rect 12124 17280 12130 17332
rect 13630 17280 13636 17332
rect 13688 17280 13694 17332
rect 14642 17280 14648 17332
rect 14700 17320 14706 17332
rect 14700 17292 14872 17320
rect 14700 17280 14706 17292
rect 10505 17255 10563 17261
rect 10505 17221 10517 17255
rect 10551 17252 10563 17255
rect 12161 17255 12219 17261
rect 10551 17224 11928 17252
rect 10551 17221 10563 17224
rect 10505 17215 10563 17221
rect 11698 17184 11704 17196
rect 10060 17156 11704 17184
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11900 17184 11928 17224
rect 12161 17221 12173 17255
rect 12207 17252 12219 17255
rect 12207 17224 13032 17252
rect 12207 17221 12219 17224
rect 12161 17215 12219 17221
rect 13004 17184 13032 17224
rect 13906 17212 13912 17264
rect 13964 17212 13970 17264
rect 14734 17212 14740 17264
rect 14792 17212 14798 17264
rect 14844 17252 14872 17292
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 15436 17292 16037 17320
rect 15436 17280 15442 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 18414 17320 18420 17332
rect 16025 17283 16083 17289
rect 16132 17292 18420 17320
rect 16132 17252 16160 17292
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 19153 17323 19211 17329
rect 19153 17289 19165 17323
rect 19199 17320 19211 17323
rect 19242 17320 19248 17332
rect 19199 17292 19248 17320
rect 19199 17289 19211 17292
rect 19153 17283 19211 17289
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 20898 17320 20904 17332
rect 19484 17292 20904 17320
rect 19484 17280 19490 17292
rect 14844 17224 16160 17252
rect 17310 17212 17316 17264
rect 17368 17252 17374 17264
rect 18138 17252 18144 17264
rect 17368 17224 18144 17252
rect 17368 17212 17374 17224
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 13924 17184 13952 17212
rect 11900 17156 12480 17184
rect 13004 17156 13952 17184
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 11054 17116 11060 17128
rect 10827 17088 11060 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10612 17048 10640 17079
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 12342 17076 12348 17128
rect 12400 17076 12406 17128
rect 12452 17116 12480 17156
rect 15102 17144 15108 17196
rect 15160 17184 15166 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15160 17156 15945 17184
rect 15160 17144 15166 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 17402 17144 17408 17196
rect 17460 17144 17466 17196
rect 19720 17193 19748 17292
rect 20898 17280 20904 17292
rect 20956 17320 20962 17332
rect 20956 17292 21312 17320
rect 20956 17280 20962 17292
rect 19978 17212 19984 17264
rect 20036 17212 20042 17264
rect 20714 17212 20720 17264
rect 20772 17212 20778 17264
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 21284 17184 21312 17292
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 21416 17292 21465 17320
rect 21416 17280 21422 17292
rect 21453 17289 21465 17292
rect 21499 17320 21511 17323
rect 21499 17292 22324 17320
rect 21499 17289 21511 17292
rect 21453 17283 21511 17289
rect 22296 17261 22324 17292
rect 22281 17255 22339 17261
rect 22281 17221 22293 17255
rect 22327 17221 22339 17255
rect 23750 17252 23756 17264
rect 23506 17238 23756 17252
rect 22281 17215 22339 17221
rect 23492 17224 23756 17238
rect 22002 17184 22008 17196
rect 21284 17156 22008 17184
rect 19705 17147 19763 17153
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 12452 17088 13308 17116
rect 12710 17048 12716 17060
rect 10612 17020 12716 17048
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 13280 17057 13308 17088
rect 13722 17076 13728 17128
rect 13780 17076 13786 17128
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 14274 17116 14280 17128
rect 13955 17088 14280 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14274 17076 14280 17088
rect 14332 17116 14338 17128
rect 14458 17116 14464 17128
rect 14332 17088 14464 17116
rect 14332 17076 14338 17088
rect 14458 17076 14464 17088
rect 14516 17076 14522 17128
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 17126 17116 17132 17128
rect 16255 17088 17132 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17116 17739 17119
rect 18414 17116 18420 17128
rect 17727 17088 18420 17116
rect 17727 17085 17739 17088
rect 17681 17079 17739 17085
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 22830 17076 22836 17128
rect 22888 17116 22894 17128
rect 23492 17116 23520 17224
rect 23750 17212 23756 17224
rect 23808 17212 23814 17264
rect 22888 17088 23520 17116
rect 22888 17076 22894 17088
rect 13265 17051 13323 17057
rect 13265 17017 13277 17051
rect 13311 17017 13323 17051
rect 13265 17011 13323 17017
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 9968 16952 11713 16980
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14829 16983 14887 16989
rect 14829 16980 14841 16983
rect 13964 16952 14841 16980
rect 13964 16940 13970 16952
rect 14829 16949 14841 16952
rect 14875 16949 14887 16983
rect 14829 16943 14887 16949
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 17770 16980 17776 16992
rect 15611 16952 17776 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 17770 16940 17776 16952
rect 17828 16940 17834 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22738 16980 22744 16992
rect 22152 16952 22744 16980
rect 22152 16940 22158 16952
rect 22738 16940 22744 16952
rect 22796 16980 22802 16992
rect 23753 16983 23811 16989
rect 23753 16980 23765 16983
rect 22796 16952 23765 16980
rect 22796 16940 22802 16952
rect 23753 16949 23765 16952
rect 23799 16949 23811 16983
rect 23753 16943 23811 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 2866 16776 2872 16788
rect 2746 16748 2872 16776
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 2746 16572 2774 16748
rect 2866 16736 2872 16748
rect 2924 16776 2930 16788
rect 9582 16776 9588 16788
rect 2924 16748 9588 16776
rect 2924 16736 2930 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 10284 16748 11100 16776
rect 10284 16736 10290 16748
rect 9125 16711 9183 16717
rect 9125 16677 9137 16711
rect 9171 16677 9183 16711
rect 9125 16671 9183 16677
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6546 16640 6552 16652
rect 5951 16612 6552 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7650 16600 7656 16652
rect 7708 16600 7714 16652
rect 2547 16544 2774 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 5626 16532 5632 16584
rect 5684 16532 5690 16584
rect 7668 16572 7696 16600
rect 9140 16584 9168 16671
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 10318 16640 10324 16652
rect 9815 16612 10324 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10778 16600 10784 16652
rect 10836 16600 10842 16652
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 11072 16640 11100 16748
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 12618 16776 12624 16788
rect 11388 16748 12624 16776
rect 11388 16736 11394 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11072 16612 11897 16640
rect 10965 16603 11023 16609
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 12161 16643 12219 16649
rect 12161 16609 12173 16643
rect 12207 16640 12219 16643
rect 12250 16640 12256 16652
rect 12207 16612 12256 16640
rect 12207 16609 12219 16612
rect 12161 16603 12219 16609
rect 7576 16544 7696 16572
rect 6178 16464 6184 16516
rect 6236 16504 6242 16516
rect 6236 16476 6394 16504
rect 6236 16464 6242 16476
rect 2590 16396 2596 16448
rect 2648 16396 2654 16448
rect 6288 16436 6316 16476
rect 6914 16436 6920 16448
rect 6288 16408 6920 16436
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7576 16436 7604 16544
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 10870 16572 10876 16584
rect 9539 16544 10876 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 10980 16572 11008 16603
rect 12250 16600 12256 16612
rect 12308 16640 12314 16652
rect 15470 16640 15476 16652
rect 12308 16612 15476 16640
rect 12308 16600 12314 16612
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 22097 16643 22155 16649
rect 22097 16609 22109 16643
rect 22143 16640 22155 16643
rect 22830 16640 22836 16652
rect 22143 16612 22836 16640
rect 22143 16609 22155 16612
rect 22097 16603 22155 16609
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 11330 16572 11336 16584
rect 10980 16544 11336 16572
rect 7653 16507 7711 16513
rect 7653 16473 7665 16507
rect 7699 16504 7711 16507
rect 10980 16504 11008 16544
rect 11330 16532 11336 16544
rect 11388 16532 11394 16584
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16572 15991 16575
rect 16206 16572 16212 16584
rect 15979 16544 16212 16572
rect 15979 16541 15991 16544
rect 15933 16535 15991 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 18322 16532 18328 16584
rect 18380 16572 18386 16584
rect 20441 16575 20499 16581
rect 20441 16572 20453 16575
rect 18380 16544 20453 16572
rect 18380 16532 18386 16544
rect 20441 16541 20453 16544
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 22649 16575 22707 16581
rect 21692 16544 22094 16572
rect 21692 16532 21698 16544
rect 7699 16476 11008 16504
rect 7699 16473 7711 16476
rect 7653 16467 7711 16473
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 11112 16476 12650 16504
rect 11112 16464 11118 16476
rect 20898 16464 20904 16516
rect 20956 16504 20962 16516
rect 21177 16507 21235 16513
rect 21177 16504 21189 16507
rect 20956 16476 21189 16504
rect 20956 16464 20962 16476
rect 21177 16473 21189 16476
rect 21223 16473 21235 16507
rect 21177 16467 21235 16473
rect 21910 16464 21916 16516
rect 21968 16464 21974 16516
rect 22066 16504 22094 16544
rect 22649 16541 22661 16575
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22664 16504 22692 16535
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 22066 16476 22692 16504
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 7576 16408 10333 16436
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 10686 16396 10692 16448
rect 10744 16396 10750 16448
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 12526 16436 12532 16448
rect 10928 16408 12532 16436
rect 10928 16396 10934 16408
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13538 16396 13544 16448
rect 13596 16436 13602 16448
rect 13633 16439 13691 16445
rect 13633 16436 13645 16439
rect 13596 16408 13645 16436
rect 13596 16396 13602 16408
rect 13633 16405 13645 16408
rect 13679 16405 13691 16439
rect 13633 16399 13691 16405
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 15749 16439 15807 16445
rect 15749 16436 15761 16439
rect 15712 16408 15761 16436
rect 15712 16396 15718 16408
rect 15749 16405 15761 16408
rect 15795 16405 15807 16439
rect 15749 16399 15807 16405
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18322 16436 18328 16448
rect 18196 16408 18328 16436
rect 18196 16396 18202 16408
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 7006 16192 7012 16244
rect 7064 16192 7070 16244
rect 7466 16192 7472 16244
rect 7524 16192 7530 16244
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 8628 16204 9137 16232
rect 8628 16192 8634 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 9217 16235 9275 16241
rect 9217 16201 9229 16235
rect 9263 16232 9275 16235
rect 9766 16232 9772 16244
rect 9263 16204 9772 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10781 16235 10839 16241
rect 10781 16201 10793 16235
rect 10827 16232 10839 16235
rect 10870 16232 10876 16244
rect 10827 16204 10876 16232
rect 10827 16201 10839 16204
rect 10781 16195 10839 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18601 16235 18659 16241
rect 18601 16232 18613 16235
rect 18472 16204 18613 16232
rect 18472 16192 18478 16204
rect 18601 16201 18613 16204
rect 18647 16201 18659 16235
rect 18601 16195 18659 16201
rect 20438 16192 20444 16244
rect 20496 16192 20502 16244
rect 21361 16235 21419 16241
rect 21361 16201 21373 16235
rect 21407 16232 21419 16235
rect 23842 16232 23848 16244
rect 21407 16204 23848 16232
rect 21407 16201 21419 16204
rect 21361 16195 21419 16201
rect 23842 16192 23848 16204
rect 23900 16192 23906 16244
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 13998 16164 14004 16176
rect 10744 16136 14004 16164
rect 10744 16124 10750 16136
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 16114 16124 16120 16176
rect 16172 16124 16178 16176
rect 17402 16164 17408 16176
rect 16868 16136 17408 16164
rect 16868 16108 16896 16136
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 20990 16124 20996 16176
rect 21048 16164 21054 16176
rect 21269 16167 21327 16173
rect 21269 16164 21281 16167
rect 21048 16136 21281 16164
rect 21048 16124 21054 16136
rect 21269 16133 21281 16136
rect 21315 16133 21327 16167
rect 21269 16127 21327 16133
rect 22281 16167 22339 16173
rect 22281 16133 22293 16167
rect 22327 16164 22339 16167
rect 22554 16164 22560 16176
rect 22327 16136 22560 16164
rect 22327 16133 22339 16136
rect 22281 16127 22339 16133
rect 22554 16124 22560 16136
rect 22612 16124 22618 16176
rect 22738 16124 22744 16176
rect 22796 16124 22802 16176
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 10873 16099 10931 16105
rect 7423 16068 8800 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 7340 16000 7573 16028
rect 7340 15988 7346 16000
rect 7561 15997 7573 16000
rect 7607 16028 7619 16031
rect 7650 16028 7656 16040
rect 7607 16000 7656 16028
rect 7607 15997 7619 16000
rect 7561 15991 7619 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 8772 15969 8800 16068
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 12802 16096 12808 16108
rect 10919 16068 12808 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15378 16096 15384 16108
rect 15243 16068 15384 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10376 16000 10977 16028
rect 10376 15988 10382 16000
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15929 8815 15963
rect 9416 15960 9444 15988
rect 12342 15960 12348 15972
rect 9416 15932 12348 15960
rect 8757 15923 8815 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 7834 15852 7840 15904
rect 7892 15892 7898 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 7892 15864 10425 15892
rect 7892 15852 7898 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 14826 15852 14832 15904
rect 14884 15852 14890 15904
rect 15212 15892 15240 16059
rect 15378 16056 15384 16068
rect 15436 16056 15442 16108
rect 16850 16056 16856 16108
rect 16908 16056 16914 16108
rect 20349 16099 20407 16105
rect 15286 15988 15292 16040
rect 15344 15988 15350 16040
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 18248 16028 18276 16082
rect 20349 16065 20361 16099
rect 20395 16096 20407 16099
rect 20806 16096 20812 16108
rect 20395 16068 20812 16096
rect 20395 16065 20407 16068
rect 20349 16059 20407 16065
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 18322 16028 18328 16040
rect 18248 16000 18328 16028
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 20530 15988 20536 16040
rect 20588 15988 20594 16040
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 22005 16031 22063 16037
rect 22005 16028 22017 16031
rect 20956 16000 22017 16028
rect 20956 15988 20962 16000
rect 22005 15997 22017 16000
rect 22051 15997 22063 16031
rect 22005 15991 22063 15997
rect 16298 15920 16304 15972
rect 16356 15920 16362 15972
rect 20346 15960 20352 15972
rect 18156 15932 20352 15960
rect 18156 15892 18184 15932
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 20438 15920 20444 15972
rect 20496 15960 20502 15972
rect 21082 15960 21088 15972
rect 20496 15932 21088 15960
rect 20496 15920 20502 15932
rect 21082 15920 21088 15932
rect 21140 15960 21146 15972
rect 21140 15932 22094 15960
rect 21140 15920 21146 15932
rect 15212 15864 18184 15892
rect 19518 15852 19524 15904
rect 19576 15852 19582 15904
rect 19981 15895 20039 15901
rect 19981 15861 19993 15895
rect 20027 15892 20039 15895
rect 21450 15892 21456 15904
rect 20027 15864 21456 15892
rect 20027 15861 20039 15864
rect 19981 15855 20039 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 22066 15892 22094 15932
rect 23753 15895 23811 15901
rect 23753 15892 23765 15895
rect 22066 15864 23765 15892
rect 23753 15861 23765 15864
rect 23799 15861 23811 15895
rect 23753 15855 23811 15861
rect 24394 15852 24400 15904
rect 24452 15852 24458 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 5776 15660 7420 15688
rect 5776 15648 5782 15660
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 6089 15555 6147 15561
rect 6089 15552 6101 15555
rect 5684 15524 6101 15552
rect 5684 15512 5690 15524
rect 6089 15521 6101 15524
rect 6135 15552 6147 15555
rect 6730 15552 6736 15564
rect 6135 15524 6736 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 7392 15552 7420 15660
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7708 15660 7849 15688
rect 7708 15648 7714 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11572 15660 11989 15688
rect 11572 15648 11578 15660
rect 11977 15657 11989 15660
rect 12023 15688 12035 15691
rect 12066 15688 12072 15700
rect 12023 15660 12072 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 22278 15688 22284 15700
rect 18187 15660 22284 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 15010 15580 15016 15632
rect 15068 15620 15074 15632
rect 18506 15620 18512 15632
rect 15068 15592 18512 15620
rect 15068 15580 15074 15592
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 19429 15623 19487 15629
rect 19429 15589 19441 15623
rect 19475 15620 19487 15623
rect 20990 15620 20996 15632
rect 19475 15592 20996 15620
rect 19475 15589 19487 15592
rect 19429 15583 19487 15589
rect 20990 15580 20996 15592
rect 21048 15580 21054 15632
rect 21453 15623 21511 15629
rect 21453 15589 21465 15623
rect 21499 15620 21511 15623
rect 23934 15620 23940 15632
rect 21499 15592 23940 15620
rect 21499 15589 21511 15592
rect 21453 15583 21511 15589
rect 23934 15580 23940 15592
rect 23992 15580 23998 15632
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 7392 15524 10517 15552
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 18414 15512 18420 15564
rect 18472 15552 18478 15564
rect 18693 15555 18751 15561
rect 18693 15552 18705 15555
rect 18472 15524 18705 15552
rect 18472 15512 18478 15524
rect 18693 15521 18705 15524
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 19886 15512 19892 15564
rect 19944 15512 19950 15564
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 20438 15552 20444 15564
rect 20119 15524 20444 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20438 15512 20444 15524
rect 20496 15512 20502 15564
rect 20809 15555 20867 15561
rect 20809 15521 20821 15555
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 14366 15444 14372 15496
rect 14424 15444 14430 15496
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 17770 15444 17776 15496
rect 17828 15484 17834 15496
rect 18601 15487 18659 15493
rect 18601 15484 18613 15487
rect 17828 15456 18613 15484
rect 17828 15444 17834 15456
rect 18601 15453 18613 15456
rect 18647 15453 18659 15487
rect 18601 15447 18659 15453
rect 20824 15428 20852 15515
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22005 15555 22063 15561
rect 21876 15524 21956 15552
rect 21876 15512 21882 15524
rect 21928 15484 21956 15524
rect 22005 15521 22017 15555
rect 22051 15552 22063 15555
rect 22094 15552 22100 15564
rect 22051 15524 22100 15552
rect 22051 15521 22063 15524
rect 22005 15515 22063 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24854 15552 24860 15564
rect 23891 15524 24860 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 22649 15487 22707 15493
rect 22649 15484 22661 15487
rect 21928 15456 22661 15484
rect 22649 15453 22661 15456
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 6365 15419 6423 15425
rect 6365 15385 6377 15419
rect 6411 15385 6423 15419
rect 6365 15379 6423 15385
rect 6380 15348 6408 15379
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 11054 15376 11060 15428
rect 11112 15376 11118 15428
rect 16945 15419 17003 15425
rect 16945 15385 16957 15419
rect 16991 15416 17003 15419
rect 17402 15416 17408 15428
rect 16991 15388 17408 15416
rect 16991 15385 17003 15388
rect 16945 15379 17003 15385
rect 17402 15376 17408 15388
rect 17460 15376 17466 15428
rect 20162 15376 20168 15428
rect 20220 15376 20226 15428
rect 20806 15376 20812 15428
rect 20864 15376 20870 15428
rect 21821 15419 21879 15425
rect 21821 15385 21833 15419
rect 21867 15416 21879 15419
rect 24394 15416 24400 15428
rect 21867 15388 24400 15416
rect 21867 15385 21879 15388
rect 21821 15379 21879 15385
rect 24394 15376 24400 15388
rect 24452 15376 24458 15428
rect 9398 15348 9404 15360
rect 6380 15320 9404 15348
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 14458 15308 14464 15360
rect 14516 15308 14522 15360
rect 18506 15308 18512 15360
rect 18564 15308 18570 15360
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 19797 15351 19855 15357
rect 19797 15348 19809 15351
rect 18932 15320 19809 15348
rect 18932 15308 18938 15320
rect 19797 15317 19809 15320
rect 19843 15317 19855 15351
rect 20180 15348 20208 15376
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 20180 15320 21925 15348
rect 19797 15311 19855 15317
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 7558 15104 7564 15156
rect 7616 15104 7622 15156
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 9122 15144 9128 15156
rect 7975 15116 9128 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9674 15144 9680 15156
rect 9416 15116 9680 15144
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 8021 15079 8079 15085
rect 8021 15076 8033 15079
rect 7892 15048 8033 15076
rect 7892 15036 7898 15048
rect 8021 15045 8033 15048
rect 8067 15045 8079 15079
rect 9416 15076 9444 15116
rect 9674 15104 9680 15116
rect 9732 15144 9738 15156
rect 10042 15144 10048 15156
rect 9732 15116 10048 15144
rect 9732 15104 9738 15116
rect 10042 15104 10048 15116
rect 10100 15144 10106 15156
rect 11054 15144 11060 15156
rect 10100 15116 11060 15144
rect 10100 15104 10106 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12860 15116 13093 15144
rect 12860 15104 12866 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 14826 15144 14832 15156
rect 13495 15116 14832 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 19058 15104 19064 15156
rect 19116 15144 19122 15156
rect 19245 15147 19303 15153
rect 19245 15144 19257 15147
rect 19116 15116 19257 15144
rect 19116 15104 19122 15116
rect 19245 15113 19257 15116
rect 19291 15113 19303 15147
rect 19245 15107 19303 15113
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19576 15116 19625 15144
rect 19576 15104 19582 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 8021 15039 8079 15045
rect 8312 15048 9522 15076
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 8312 15008 8340 15048
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 13541 15079 13599 15085
rect 13541 15045 13553 15079
rect 13587 15076 13599 15079
rect 13630 15076 13636 15088
rect 13587 15048 13636 15076
rect 13587 15045 13599 15048
rect 13541 15039 13599 15045
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 15286 15036 15292 15088
rect 15344 15076 15350 15088
rect 15838 15076 15844 15088
rect 15344 15048 15844 15076
rect 15344 15036 15350 15048
rect 15838 15036 15844 15048
rect 15896 15076 15902 15088
rect 19705 15079 19763 15085
rect 19705 15076 19717 15079
rect 15896 15048 19717 15076
rect 15896 15036 15902 15048
rect 19705 15045 19717 15048
rect 19751 15045 19763 15079
rect 19705 15039 19763 15045
rect 23293 15079 23351 15085
rect 23293 15045 23305 15079
rect 23339 15076 23351 15079
rect 24854 15076 24860 15088
rect 23339 15048 24860 15076
rect 23339 15045 23351 15048
rect 23293 15039 23351 15045
rect 24854 15036 24860 15048
rect 24912 15036 24918 15088
rect 13354 15008 13360 15020
rect 6972 14980 8340 15008
rect 12728 14980 13360 15008
rect 6972 14968 6978 14980
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14940 8263 14943
rect 8570 14940 8576 14952
rect 8251 14912 8576 14940
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 8754 14900 8760 14952
rect 8812 14900 8818 14952
rect 9030 14900 9036 14952
rect 9088 14900 9094 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 12621 14943 12679 14949
rect 12621 14940 12633 14943
rect 9824 14912 12633 14940
rect 9824 14900 9830 14912
rect 12621 14909 12633 14912
rect 12667 14909 12679 14943
rect 12621 14903 12679 14909
rect 12434 14832 12440 14884
rect 12492 14872 12498 14884
rect 12728 14872 12756 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 13504 14980 17417 15008
rect 13504 14968 13510 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18564 14980 18797 15008
rect 18564 14968 18570 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 15008 21051 15011
rect 21174 15008 21180 15020
rect 21039 14980 21180 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 21174 14968 21180 14980
rect 21232 14968 21238 15020
rect 22186 14968 22192 15020
rect 22244 14968 22250 15020
rect 24121 15011 24179 15017
rect 24121 14977 24133 15011
rect 24167 15008 24179 15011
rect 24210 15008 24216 15020
rect 24167 14980 24216 15008
rect 24167 14977 24179 14980
rect 24121 14971 24179 14977
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 13538 14940 13544 14952
rect 12860 14912 13544 14940
rect 12860 14900 12866 14912
rect 13538 14900 13544 14912
rect 13596 14940 13602 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13596 14912 13645 14940
rect 13596 14900 13602 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 17497 14943 17555 14949
rect 17497 14940 17509 14943
rect 14148 14912 17509 14940
rect 14148 14900 14154 14912
rect 17497 14909 17509 14912
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 17589 14943 17647 14949
rect 17589 14909 17601 14943
rect 17635 14909 17647 14943
rect 17589 14903 17647 14909
rect 19889 14943 19947 14949
rect 19889 14909 19901 14943
rect 19935 14940 19947 14943
rect 22462 14940 22468 14952
rect 19935 14912 22468 14940
rect 19935 14909 19947 14912
rect 19889 14903 19947 14909
rect 12492 14844 12756 14872
rect 12492 14832 12498 14844
rect 13262 14832 13268 14884
rect 13320 14872 13326 14884
rect 13320 14844 13584 14872
rect 13320 14832 13326 14844
rect 13556 14816 13584 14844
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17604 14872 17632 14903
rect 22462 14900 22468 14912
rect 22520 14900 22526 14952
rect 24762 14900 24768 14952
rect 24820 14900 24826 14952
rect 17276 14844 17632 14872
rect 17276 14832 17282 14844
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 10376 14776 10517 14804
rect 10376 14764 10382 14776
rect 10505 14773 10517 14776
rect 10551 14773 10563 14807
rect 10505 14767 10563 14773
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 13354 14804 13360 14816
rect 11480 14776 13360 14804
rect 11480 14764 11486 14776
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 13538 14764 13544 14816
rect 13596 14764 13602 14816
rect 17037 14807 17095 14813
rect 17037 14773 17049 14807
rect 17083 14804 17095 14807
rect 18322 14804 18328 14816
rect 17083 14776 18328 14804
rect 17083 14773 17095 14776
rect 17037 14767 17095 14773
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 20806 14764 20812 14816
rect 20864 14764 20870 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 9217 14603 9275 14609
rect 9217 14569 9229 14603
rect 9263 14600 9275 14603
rect 9582 14600 9588 14612
rect 9263 14572 9588 14600
rect 9263 14569 9275 14572
rect 9217 14563 9275 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10670 14603 10728 14609
rect 10670 14600 10682 14603
rect 10560 14572 10682 14600
rect 10560 14560 10566 14572
rect 10670 14569 10682 14572
rect 10716 14569 10728 14603
rect 10670 14563 10728 14569
rect 11790 14560 11796 14612
rect 11848 14600 11854 14612
rect 12805 14603 12863 14609
rect 12805 14600 12817 14603
rect 11848 14572 12817 14600
rect 11848 14560 11854 14572
rect 12805 14569 12817 14572
rect 12851 14569 12863 14603
rect 12805 14563 12863 14569
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 17126 14600 17132 14612
rect 16807 14572 17132 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 12676 14504 13400 14532
rect 12676 14492 12682 14504
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 8754 14464 8760 14476
rect 6871 14436 8760 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9088 14436 9873 14464
rect 9088 14424 9094 14436
rect 9861 14433 9873 14436
rect 9907 14464 9919 14467
rect 12802 14464 12808 14476
rect 9907 14436 12808 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 13372 14473 13400 14504
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14332 14436 15025 14464
rect 14332 14424 14338 14436
rect 15013 14433 15025 14436
rect 15059 14464 15071 14467
rect 16850 14464 16856 14476
rect 15059 14436 16856 14464
rect 15059 14433 15071 14436
rect 15013 14427 15071 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 8772 14396 8800 14424
rect 9398 14396 9404 14408
rect 8772 14368 9404 14396
rect 9398 14356 9404 14368
rect 9456 14396 9462 14408
rect 10226 14396 10232 14408
rect 9456 14368 10232 14396
rect 9456 14356 9462 14368
rect 10226 14356 10232 14368
rect 10284 14396 10290 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10284 14368 10425 14396
rect 10284 14356 10290 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13136 14368 13185 14396
rect 13136 14356 13142 14368
rect 13173 14365 13185 14368
rect 13219 14396 13231 14399
rect 13906 14396 13912 14408
rect 13219 14368 13912 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13906 14356 13912 14368
rect 13964 14396 13970 14408
rect 14826 14396 14832 14408
rect 13964 14368 14832 14396
rect 13964 14356 13970 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 18598 14396 18604 14408
rect 17543 14368 18604 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 20622 14356 20628 14408
rect 20680 14356 20686 14408
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 22428 14368 23397 14396
rect 22428 14356 22434 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 7101 14331 7159 14337
rect 7101 14297 7113 14331
rect 7147 14297 7159 14331
rect 7101 14291 7159 14297
rect 7116 14260 7144 14291
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 7558 14328 7564 14340
rect 7248 14300 7564 14328
rect 7248 14288 7254 14300
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 10318 14328 10324 14340
rect 8496 14300 10324 14328
rect 8496 14260 8524 14300
rect 10318 14288 10324 14300
rect 10376 14288 10382 14340
rect 11146 14288 11152 14340
rect 11204 14288 11210 14340
rect 13265 14331 13323 14337
rect 13265 14297 13277 14331
rect 13311 14328 13323 14331
rect 13446 14328 13452 14340
rect 13311 14300 13452 14328
rect 13311 14297 13323 14300
rect 13265 14291 13323 14297
rect 13446 14288 13452 14300
rect 13504 14288 13510 14340
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 16022 14288 16028 14340
rect 16080 14288 16086 14340
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18049 14331 18107 14337
rect 18049 14328 18061 14331
rect 18012 14300 18061 14328
rect 18012 14288 18018 14300
rect 18049 14297 18061 14300
rect 18095 14297 18107 14331
rect 18049 14291 18107 14297
rect 18233 14331 18291 14337
rect 18233 14297 18245 14331
rect 18279 14328 18291 14331
rect 21266 14328 21272 14340
rect 18279 14300 21272 14328
rect 18279 14297 18291 14300
rect 18233 14291 18291 14297
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 7116 14232 8524 14260
rect 8570 14220 8576 14272
rect 8628 14220 8634 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9585 14263 9643 14269
rect 9585 14260 9597 14263
rect 9088 14232 9597 14260
rect 9088 14220 9094 14232
rect 9585 14229 9597 14232
rect 9631 14229 9643 14263
rect 9585 14223 9643 14229
rect 9674 14220 9680 14272
rect 9732 14220 9738 14272
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14260 12219 14263
rect 12342 14260 12348 14272
rect 12207 14232 12348 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 17313 14263 17371 14269
rect 17313 14229 17325 14263
rect 17359 14260 17371 14263
rect 17402 14260 17408 14272
rect 17359 14232 17408 14260
rect 17359 14229 17371 14232
rect 17313 14223 17371 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20441 14263 20499 14269
rect 20441 14260 20453 14263
rect 20128 14232 20453 14260
rect 20128 14220 20134 14232
rect 20441 14229 20453 14232
rect 20487 14229 20499 14263
rect 20441 14223 20499 14229
rect 23201 14263 23259 14269
rect 23201 14229 23213 14263
rect 23247 14260 23259 14263
rect 23382 14260 23388 14272
rect 23247 14232 23388 14260
rect 23247 14229 23259 14232
rect 23201 14223 23259 14229
rect 23382 14220 23388 14232
rect 23440 14220 23446 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9490 14056 9496 14068
rect 9272 14028 9496 14056
rect 9272 14016 9278 14028
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 13078 14016 13084 14068
rect 13136 14016 13142 14068
rect 13173 14059 13231 14065
rect 13173 14025 13185 14059
rect 13219 14056 13231 14059
rect 13446 14056 13452 14068
rect 13219 14028 13452 14056
rect 13219 14025 13231 14028
rect 13173 14019 13231 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 17310 14056 17316 14068
rect 13955 14028 17316 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18414 14056 18420 14068
rect 17512 14028 18420 14056
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 9125 13991 9183 13997
rect 9125 13988 9137 13991
rect 8628 13960 9137 13988
rect 8628 13948 8634 13960
rect 9125 13957 9137 13960
rect 9171 13957 9183 13991
rect 9125 13951 9183 13957
rect 10134 13948 10140 14000
rect 10192 13948 10198 14000
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 10836 13960 14289 13988
rect 10836 13948 10842 13960
rect 14277 13957 14289 13960
rect 14323 13957 14335 13991
rect 14277 13951 14335 13957
rect 15289 13991 15347 13997
rect 15289 13957 15301 13991
rect 15335 13988 15347 13991
rect 15562 13988 15568 14000
rect 15335 13960 15568 13988
rect 15335 13957 15347 13960
rect 15289 13951 15347 13957
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 16022 13988 16028 14000
rect 15712 13960 16028 13988
rect 15712 13948 15718 13960
rect 16022 13948 16028 13960
rect 16080 13988 16086 14000
rect 17512 13988 17540 14028
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18690 14056 18696 14068
rect 18647 14028 18696 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 21048 14028 21189 14056
rect 21048 14016 21054 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 22005 14059 22063 14065
rect 22005 14025 22017 14059
rect 22051 14056 22063 14059
rect 24578 14056 24584 14068
rect 22051 14028 24584 14056
rect 22051 14025 22063 14028
rect 22005 14019 22063 14025
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 16080 13960 17618 13988
rect 16080 13948 16086 13960
rect 19794 13948 19800 14000
rect 19852 13988 19858 14000
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 19852 13960 19901 13988
rect 19852 13948 19858 13960
rect 19889 13957 19901 13960
rect 19935 13957 19947 13991
rect 19889 13951 19947 13957
rect 21085 13991 21143 13997
rect 21085 13957 21097 13991
rect 21131 13988 21143 13991
rect 23290 13988 23296 14000
rect 21131 13960 23296 13988
rect 21131 13957 21143 13960
rect 21085 13951 21143 13957
rect 23290 13948 23296 13960
rect 23348 13948 23354 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 2590 13920 2596 13932
rect 1811 13892 2596 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8812 13892 8861 13920
rect 8812 13880 8818 13892
rect 8849 13889 8861 13892
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10870 13920 10876 13932
rect 10560 13892 10876 13920
rect 10560 13880 10566 13892
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 13446 13920 13452 13932
rect 12032 13892 13452 13920
rect 12032 13880 12038 13892
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 14148 13892 14381 13920
rect 14148 13880 14154 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 16850 13880 16856 13932
rect 16908 13880 16914 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18782 13920 18788 13932
rect 18472 13892 18788 13920
rect 18472 13880 18478 13892
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 21542 13920 21548 13932
rect 20119 13892 21548 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 22278 13920 22284 13932
rect 22235 13892 22284 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12768 13824 13277 13852
rect 12768 13812 12774 13824
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13265 13815 13323 13821
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 15473 13855 15531 13861
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 16666 13852 16672 13864
rect 15519 13824 16672 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 13280 13784 13308 13815
rect 14366 13784 14372 13796
rect 13280 13756 14372 13784
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 14568 13728 14596 13815
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 20254 13744 20260 13796
rect 20312 13784 20318 13796
rect 21284 13784 21312 13815
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22848 13852 22876 13883
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23532 13892 23949 13920
rect 23532 13880 23538 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 21508 13824 22876 13852
rect 21508 13812 21514 13824
rect 20312 13756 21312 13784
rect 20312 13744 20318 13756
rect 14550 13676 14556 13728
rect 14608 13676 14614 13728
rect 18782 13676 18788 13728
rect 18840 13716 18846 13728
rect 19245 13719 19303 13725
rect 19245 13716 19257 13719
rect 18840 13688 19257 13716
rect 18840 13676 18846 13688
rect 19245 13685 19257 13688
rect 19291 13685 19303 13719
rect 19245 13679 19303 13685
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 21450 13716 21456 13728
rect 21324 13688 21456 13716
rect 21324 13676 21330 13688
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 22646 13676 22652 13728
rect 22704 13676 22710 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13538 13512 13544 13524
rect 13320 13484 13544 13512
rect 13320 13472 13326 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 21266 13512 21272 13524
rect 18187 13484 21272 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 23290 13472 23296 13524
rect 23348 13472 23354 13524
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 13446 13444 13452 13456
rect 12023 13416 13452 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 18874 13444 18880 13456
rect 16080 13416 18880 13444
rect 16080 13404 16086 13416
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7742 13376 7748 13388
rect 7156 13348 7748 13376
rect 7156 13336 7162 13348
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 11204 13348 12541 13376
rect 11204 13336 11210 13348
rect 12529 13345 12541 13348
rect 12575 13345 12587 13379
rect 12529 13339 12587 13345
rect 18322 13336 18328 13388
rect 18380 13376 18386 13388
rect 18601 13379 18659 13385
rect 18601 13376 18613 13379
rect 18380 13348 18613 13376
rect 18380 13336 18386 13348
rect 18601 13345 18613 13348
rect 18647 13345 18659 13379
rect 18601 13339 18659 13345
rect 18690 13336 18696 13388
rect 18748 13336 18754 13388
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21634 13376 21640 13388
rect 20680 13348 21640 13376
rect 20680 13336 20686 13348
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 9088 13280 12357 13308
rect 9088 13268 9094 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13308 12495 13311
rect 13814 13308 13820 13320
rect 12483 13280 13820 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 14918 13268 14924 13320
rect 14976 13268 14982 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13308 16911 13311
rect 17218 13308 17224 13320
rect 16899 13280 17224 13308
rect 16899 13277 16911 13280
rect 16853 13271 16911 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 18782 13308 18788 13320
rect 18555 13280 18788 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 19242 13268 19248 13320
rect 19300 13308 19306 13320
rect 20898 13308 20904 13320
rect 19300 13280 20904 13308
rect 19300 13268 19306 13280
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 7558 13200 7564 13252
rect 7616 13200 7622 13252
rect 8573 13175 8631 13181
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 9674 13172 9680 13184
rect 8619 13144 9680 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 13832 13172 13860 13268
rect 15105 13243 15163 13249
rect 15105 13209 15117 13243
rect 15151 13240 15163 13243
rect 16114 13240 16120 13252
rect 15151 13212 16120 13240
rect 15151 13209 15163 13212
rect 15105 13203 15163 13209
rect 16114 13200 16120 13212
rect 16172 13200 16178 13252
rect 19610 13200 19616 13252
rect 19668 13240 19674 13252
rect 19705 13243 19763 13249
rect 19705 13240 19717 13243
rect 19668 13212 19717 13240
rect 19668 13200 19674 13212
rect 19705 13209 19717 13212
rect 19751 13209 19763 13243
rect 19705 13203 19763 13209
rect 19889 13243 19947 13249
rect 19889 13209 19901 13243
rect 19935 13240 19947 13243
rect 20530 13240 20536 13252
rect 19935 13212 20536 13240
rect 19935 13209 19947 13212
rect 19889 13203 19947 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 21082 13200 21088 13252
rect 21140 13240 21146 13252
rect 21177 13243 21235 13249
rect 21177 13240 21189 13243
rect 21140 13212 21189 13240
rect 21140 13200 21146 13212
rect 21177 13209 21189 13212
rect 21223 13209 21235 13243
rect 21177 13203 21235 13209
rect 21634 13200 21640 13252
rect 21692 13200 21698 13252
rect 18506 13172 18512 13184
rect 13832 13144 18512 13172
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 22649 13175 22707 13181
rect 22649 13172 22661 13175
rect 20312 13144 22661 13172
rect 20312 13132 20318 13144
rect 22649 13141 22661 13144
rect 22695 13141 22707 13175
rect 22649 13135 22707 13141
rect 23750 13132 23756 13184
rect 23808 13132 23814 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9401 12971 9459 12977
rect 9401 12968 9413 12971
rect 9364 12940 9413 12968
rect 9364 12928 9370 12940
rect 9401 12937 9413 12940
rect 9447 12937 9459 12971
rect 9401 12931 9459 12937
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11756 12940 11805 12968
rect 11756 12928 11762 12940
rect 11793 12937 11805 12940
rect 11839 12937 11851 12971
rect 11793 12931 11851 12937
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15344 12940 16037 12968
rect 15344 12928 15350 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 12253 12903 12311 12909
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 12802 12900 12808 12912
rect 12299 12872 12808 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 13633 12903 13691 12909
rect 13633 12900 13645 12903
rect 13412 12872 13645 12900
rect 13412 12860 13418 12872
rect 13633 12869 13645 12872
rect 13679 12869 13691 12903
rect 13633 12863 13691 12869
rect 14550 12860 14556 12912
rect 14608 12860 14614 12912
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 6604 12804 9321 12832
rect 6604 12792 6610 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 13538 12832 13544 12844
rect 12207 12804 13544 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 9674 12764 9680 12776
rect 9631 12736 9680 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 16040 12764 16068 12931
rect 17218 12928 17224 12980
rect 17276 12928 17282 12980
rect 17310 12928 17316 12980
rect 17368 12928 17374 12980
rect 18506 12928 18512 12980
rect 18564 12928 18570 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 19168 12940 21465 12968
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 18380 12872 18736 12900
rect 18380 12860 18386 12872
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 16264 12804 18429 12832
rect 16264 12792 16270 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 18708 12773 18736 12872
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16040 12736 17417 12764
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 18693 12767 18751 12773
rect 18693 12733 18705 12767
rect 18739 12764 18751 12767
rect 19168 12764 19196 12940
rect 21453 12937 21465 12940
rect 21499 12937 21511 12971
rect 21453 12931 21511 12937
rect 19981 12903 20039 12909
rect 19981 12869 19993 12903
rect 20027 12900 20039 12903
rect 20254 12900 20260 12912
rect 20027 12872 20260 12900
rect 20027 12869 20039 12872
rect 19981 12863 20039 12869
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 20622 12860 20628 12912
rect 20680 12860 20686 12912
rect 23293 12903 23351 12909
rect 23293 12869 23305 12903
rect 23339 12900 23351 12903
rect 24854 12900 24860 12912
rect 23339 12872 24860 12900
rect 23339 12869 23351 12872
rect 23293 12863 23351 12869
rect 24854 12860 24860 12872
rect 24912 12860 24918 12912
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 22888 12804 23949 12832
rect 22888 12792 22894 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 18739 12736 19196 12764
rect 18739 12733 18751 12736
rect 18693 12727 18751 12733
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19300 12736 19717 12764
rect 19300 12724 19306 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 13817 12699 13875 12705
rect 13817 12665 13829 12699
rect 13863 12696 13875 12699
rect 14274 12696 14280 12708
rect 13863 12668 14280 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 19518 12696 19524 12708
rect 16899 12668 19524 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12628 8999 12631
rect 10962 12628 10968 12640
rect 8987 12600 10968 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12628 18107 12631
rect 19702 12628 19708 12640
rect 18095 12600 19708 12628
rect 18095 12597 18107 12600
rect 18049 12591 18107 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 11146 12384 11152 12436
rect 11204 12384 11210 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 14918 12424 14924 12436
rect 13688 12396 14924 12424
rect 13688 12384 13694 12396
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16482 12384 16488 12436
rect 16540 12424 16546 12436
rect 16574 12424 16580 12436
rect 16540 12396 16580 12424
rect 16540 12384 16546 12396
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 20901 12427 20959 12433
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 22094 12424 22100 12436
rect 20947 12396 22100 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 4890 12356 4896 12368
rect 2832 12328 4896 12356
rect 2832 12316 2838 12328
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 14734 12356 14740 12368
rect 13504 12328 14740 12356
rect 13504 12316 13510 12328
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 16209 12359 16267 12365
rect 16209 12325 16221 12359
rect 16255 12325 16267 12359
rect 16209 12319 16267 12325
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11020 12260 13768 12288
rect 11020 12248 11026 12260
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 11940 12192 12817 12220
rect 11940 12180 11946 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13630 12220 13636 12232
rect 13035 12192 13636 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 13740 12220 13768 12260
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 13872 12260 14841 12288
rect 13872 12248 13878 12260
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 16224 12288 16252 12319
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 20070 12356 20076 12368
rect 16448 12328 20076 12356
rect 16448 12316 16454 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 16224 12260 16574 12288
rect 14829 12251 14887 12257
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 13740 12192 16405 12220
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16546 12220 16574 12260
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 20622 12288 20628 12300
rect 19392 12260 20628 12288
rect 19392 12248 19398 12260
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 16546 12192 21097 12220
rect 16393 12183 16451 12189
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 22370 12180 22376 12232
rect 22428 12220 22434 12232
rect 22649 12223 22707 12229
rect 22649 12220 22661 12223
rect 22428 12192 22661 12220
rect 22428 12180 22434 12192
rect 22649 12189 22661 12192
rect 22695 12189 22707 12223
rect 22649 12183 22707 12189
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24636 12192 24777 12220
rect 24636 12180 24642 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 10134 12112 10140 12164
rect 10192 12112 10198 12164
rect 13354 12112 13360 12164
rect 13412 12152 13418 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13412 12124 13553 12152
rect 13412 12112 13418 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 14734 12112 14740 12164
rect 14792 12112 14798 12164
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15565 12155 15623 12161
rect 15565 12152 15577 12155
rect 15252 12124 15577 12152
rect 15252 12112 15258 12124
rect 15565 12121 15577 12124
rect 15611 12121 15623 12155
rect 15565 12115 15623 12121
rect 15749 12155 15807 12161
rect 15749 12121 15761 12155
rect 15795 12152 15807 12155
rect 16758 12152 16764 12164
rect 15795 12124 16764 12152
rect 15795 12121 15807 12124
rect 15749 12115 15807 12121
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 17957 12155 18015 12161
rect 17957 12121 17969 12155
rect 18003 12121 18015 12155
rect 17957 12115 18015 12121
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18690 12152 18696 12164
rect 18187 12124 18696 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 12492 12056 13645 12084
rect 12492 12044 12498 12056
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 14277 12087 14335 12093
rect 14277 12053 14289 12087
rect 14323 12084 14335 12087
rect 14366 12084 14372 12096
rect 14323 12056 14372 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14642 12044 14648 12096
rect 14700 12044 14706 12096
rect 17972 12084 18000 12115
rect 18690 12112 18696 12124
rect 18748 12112 18754 12164
rect 19426 12112 19432 12164
rect 19484 12152 19490 12164
rect 19521 12155 19579 12161
rect 19521 12152 19533 12155
rect 19484 12124 19533 12152
rect 19484 12112 19490 12124
rect 19521 12121 19533 12124
rect 19567 12121 19579 12155
rect 19521 12115 19579 12121
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 25314 12152 25320 12164
rect 23891 12124 25320 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 25314 12112 25320 12124
rect 25372 12112 25378 12164
rect 18414 12084 18420 12096
rect 17972 12056 18420 12084
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19610 12044 19616 12096
rect 19668 12044 19674 12096
rect 24578 12044 24584 12096
rect 24636 12044 24642 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13814 11880 13820 11892
rect 12912 11852 13820 11880
rect 12912 11821 12940 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14550 11880 14556 11892
rect 14415 11852 14556 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14918 11840 14924 11892
rect 14976 11840 14982 11892
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15335 11852 17080 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 12897 11815 12955 11821
rect 12897 11781 12909 11815
rect 12943 11781 12955 11815
rect 15654 11812 15660 11824
rect 12897 11775 12955 11781
rect 14568 11784 15660 11812
rect 14568 11744 14596 11784
rect 15654 11772 15660 11784
rect 15712 11812 15718 11824
rect 17052 11812 17080 11852
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 17184 11852 18981 11880
rect 17184 11840 17190 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 18969 11843 19027 11849
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11849 19671 11883
rect 19613 11843 19671 11849
rect 17402 11812 17408 11824
rect 15712 11784 16620 11812
rect 17052 11784 17408 11812
rect 15712 11772 15718 11784
rect 14030 11730 14596 11744
rect 14016 11716 14596 11730
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 11238 11676 11244 11688
rect 9456 11648 11244 11676
rect 9456 11636 9462 11648
rect 11238 11636 11244 11648
rect 11296 11676 11302 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 11296 11648 12633 11676
rect 11296 11636 11302 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 14016 11676 14044 11716
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 14700 11716 16313 11744
rect 14700 11704 14706 11716
rect 16301 11713 16313 11716
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 12621 11639 12679 11645
rect 12728 11648 14044 11676
rect 11974 11568 11980 11620
rect 12032 11608 12038 11620
rect 12728 11608 12756 11648
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15344 11648 15393 11676
rect 15344 11636 15350 11648
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 12032 11580 12756 11608
rect 15396 11608 15424 11639
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 16206 11608 16212 11620
rect 15396 11580 16212 11608
rect 12032 11568 12038 11580
rect 16206 11568 16212 11580
rect 16264 11568 16270 11620
rect 16592 11540 16620 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 19334 11812 19340 11824
rect 18722 11784 19340 11812
rect 19334 11772 19340 11784
rect 19392 11772 19398 11824
rect 19628 11812 19656 11843
rect 22370 11840 22376 11892
rect 22428 11840 22434 11892
rect 19628 11784 23428 11812
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16908 11716 17233 11744
rect 16908 11704 16914 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19576 11716 19809 11744
rect 19576 11704 19582 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 20346 11704 20352 11756
rect 20404 11704 20410 11756
rect 22554 11704 22560 11756
rect 22612 11704 22618 11756
rect 23400 11753 23428 11784
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11713 23443 11747
rect 23385 11707 23443 11713
rect 23842 11704 23848 11756
rect 23900 11744 23906 11756
rect 23937 11747 23995 11753
rect 23937 11744 23949 11747
rect 23900 11716 23949 11744
rect 23900 11704 23906 11716
rect 23937 11713 23949 11716
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11676 17555 11679
rect 19978 11676 19984 11688
rect 17543 11648 19984 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 24670 11636 24676 11688
rect 24728 11636 24734 11688
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19794 11608 19800 11620
rect 19392 11580 19800 11608
rect 19392 11568 19398 11580
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 20533 11611 20591 11617
rect 20533 11577 20545 11611
rect 20579 11608 20591 11611
rect 22830 11608 22836 11620
rect 20579 11580 22836 11608
rect 20579 11577 20591 11580
rect 20533 11571 20591 11577
rect 22830 11568 22836 11580
rect 22888 11568 22894 11620
rect 19426 11540 19432 11552
rect 16592 11512 19432 11540
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 23201 11543 23259 11549
rect 23201 11509 23213 11543
rect 23247 11540 23259 11543
rect 23934 11540 23940 11552
rect 23247 11512 23940 11540
rect 23247 11509 23259 11512
rect 23201 11503 23259 11509
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13814 11336 13820 11348
rect 13035 11308 13820 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 22554 11336 22560 11348
rect 18187 11308 22560 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 23290 11296 23296 11348
rect 23348 11336 23354 11348
rect 24765 11339 24823 11345
rect 24765 11336 24777 11339
rect 23348 11308 24777 11336
rect 23348 11296 23354 11308
rect 24765 11305 24777 11308
rect 24811 11305 24823 11339
rect 24765 11299 24823 11305
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 10928 11240 11376 11268
rect 10928 11228 10934 11240
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11348 11200 11376 11240
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 14277 11271 14335 11277
rect 14277 11268 14289 11271
rect 13596 11240 14289 11268
rect 13596 11228 13602 11240
rect 14277 11237 14289 11240
rect 14323 11237 14335 11271
rect 14277 11231 14335 11237
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 19429 11271 19487 11277
rect 14424 11240 16574 11268
rect 14424 11228 14430 11240
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 11348 11172 14933 11200
rect 14921 11169 14933 11172
rect 14967 11200 14979 11203
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 14967 11172 16037 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11132 14703 11135
rect 15746 11132 15752 11144
rect 14691 11104 15752 11132
rect 14691 11101 14703 11104
rect 14645 11095 14703 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16390 11132 16396 11144
rect 15887 11104 16396 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16546 11132 16574 11240
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 22186 11268 22192 11280
rect 19475 11240 22192 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 19760 11172 19901 11200
rect 19760 11160 19766 11172
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20714 11160 20720 11212
rect 20772 11200 20778 11212
rect 20772 11172 21864 11200
rect 20772 11160 20778 11172
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 16546 11104 18337 11132
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20809 11135 20867 11141
rect 20809 11132 20821 11135
rect 19843 11104 20821 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 20809 11101 20821 11104
rect 20855 11101 20867 11135
rect 21836 11132 21864 11172
rect 22646 11160 22652 11212
rect 22704 11200 22710 11212
rect 22704 11172 24072 11200
rect 22704 11160 22710 11172
rect 24044 11141 24072 11172
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 21836 11104 22937 11132
rect 20809 11095 20867 11101
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 24029 11135 24087 11141
rect 24029 11101 24041 11135
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 10192 11036 11100 11064
rect 10192 11024 10198 11036
rect 11072 10996 11100 11036
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11517 11067 11575 11073
rect 11517 11064 11529 11067
rect 11204 11036 11529 11064
rect 11204 11024 11210 11036
rect 11517 11033 11529 11036
rect 11563 11033 11575 11067
rect 11974 11064 11980 11076
rect 11517 11027 11575 11033
rect 11624 11036 11980 11064
rect 11624 10996 11652 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 12802 11024 12808 11076
rect 12860 11064 12866 11076
rect 15933 11067 15991 11073
rect 12860 11036 15516 11064
rect 12860 11024 12866 11036
rect 11072 10968 11652 10996
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 15010 10996 15016 11008
rect 14792 10968 15016 10996
rect 14792 10956 14798 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15488 11005 15516 11036
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16022 11064 16028 11076
rect 15979 11036 16028 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 23382 11024 23388 11076
rect 23440 11064 23446 11076
rect 24673 11067 24731 11073
rect 24673 11064 24685 11067
rect 23440 11036 24685 11064
rect 23440 11024 23446 11036
rect 24673 11033 24685 11036
rect 24719 11033 24731 11067
rect 24673 11027 24731 11033
rect 15473 10999 15531 11005
rect 15473 10965 15485 10999
rect 15519 10965 15531 10999
rect 15473 10959 15531 10965
rect 22738 10956 22744 11008
rect 22796 10956 22802 11008
rect 23842 10956 23848 11008
rect 23900 10956 23906 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 19242 10792 19248 10804
rect 18064 10764 19248 10792
rect 18064 10665 18092 10764
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19797 10795 19855 10801
rect 19797 10761 19809 10795
rect 19843 10792 19855 10795
rect 19978 10792 19984 10804
rect 19843 10764 19984 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 18322 10684 18328 10736
rect 18380 10684 18386 10736
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19794 10656 19800 10668
rect 19484 10628 19800 10656
rect 19484 10616 19490 10628
rect 19794 10616 19800 10628
rect 19852 10616 19858 10668
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 21085 10455 21143 10461
rect 21085 10421 21097 10455
rect 21131 10452 21143 10455
rect 24670 10452 24676 10464
rect 21131 10424 24676 10452
rect 21131 10421 21143 10424
rect 21085 10415 21143 10421
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 23808 10084 24808 10112
rect 23808 10072 23814 10084
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 9916 10016 11621 10044
rect 9916 10004 9922 10016
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10044 17003 10047
rect 20162 10044 20168 10056
rect 16991 10016 20168 10044
rect 16991 10013 17003 10016
rect 16945 10007 17003 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10044 22891 10047
rect 24578 10044 24584 10056
rect 22879 10016 24584 10044
rect 22879 10013 22891 10016
rect 22833 10007 22891 10013
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 24780 10053 24808 10084
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 23845 9979 23903 9985
rect 23845 9945 23857 9979
rect 23891 9976 23903 9979
rect 24946 9976 24952 9988
rect 23891 9948 24952 9976
rect 23891 9945 23903 9948
rect 23845 9939 23903 9945
rect 24946 9936 24952 9948
rect 25004 9936 25010 9988
rect 11698 9868 11704 9920
rect 11756 9868 11762 9920
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 17037 9911 17095 9917
rect 17037 9908 17049 9911
rect 14884 9880 17049 9908
rect 14884 9868 14890 9880
rect 17037 9877 17049 9880
rect 17083 9877 17095 9911
rect 17037 9871 17095 9877
rect 24578 9868 24584 9920
rect 24636 9868 24642 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14277 9639 14335 9645
rect 14277 9636 14289 9639
rect 14240 9608 14289 9636
rect 14240 9596 14246 9608
rect 14277 9605 14289 9608
rect 14323 9605 14335 9639
rect 14277 9599 14335 9605
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9568 6055 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6043 9540 6929 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23624 9540 23949 9568
rect 23624 9528 23630 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 5592 9472 7021 9500
rect 5592 9460 5598 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 6546 9392 6552 9444
rect 6604 9392 6610 9444
rect 14461 9435 14519 9441
rect 14461 9401 14473 9435
rect 14507 9432 14519 9435
rect 15194 9432 15200 9444
rect 14507 9404 15200 9432
rect 14507 9401 14519 9404
rect 14461 9395 14519 9401
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9364 22063 9367
rect 24026 9364 24032 9376
rect 22051 9336 24032 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 5902 9160 5908 9172
rect 3108 9132 5908 9160
rect 3108 9120 3114 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 22738 8984 22744 9036
rect 22796 9024 22802 9036
rect 22796 8996 24808 9024
rect 22796 8984 22802 8996
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15988 8928 16129 8956
rect 15988 8916 15994 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8956 18567 8959
rect 18782 8956 18788 8968
rect 18555 8928 18788 8956
rect 18555 8925 18567 8928
rect 18509 8919 18567 8925
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 24026 8916 24032 8968
rect 24084 8916 24090 8968
rect 24780 8965 24808 8996
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 17770 8888 17776 8900
rect 16347 8860 17776 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 17770 8848 17776 8860
rect 17828 8848 17834 8900
rect 18693 8891 18751 8897
rect 18693 8857 18705 8891
rect 18739 8888 18751 8891
rect 20714 8888 20720 8900
rect 18739 8860 20720 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 7558 8820 7564 8832
rect 5868 8792 7564 8820
rect 5868 8780 5874 8792
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 22830 8780 22836 8832
rect 22888 8820 22894 8832
rect 23845 8823 23903 8829
rect 23845 8820 23857 8823
rect 22888 8792 23857 8820
rect 22888 8780 22894 8792
rect 23845 8789 23857 8792
rect 23891 8789 23903 8823
rect 23845 8783 23903 8789
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 24176 8792 24593 8820
rect 24176 8780 24182 8792
rect 24581 8789 24593 8792
rect 24627 8789 24639 8823
rect 24581 8783 24639 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 6822 8616 6828 8628
rect 3896 8588 6828 8616
rect 3896 8489 3924 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16022 8616 16028 8628
rect 15804 8588 16028 8616
rect 15804 8576 15810 8588
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 5810 8548 5816 8560
rect 5382 8520 5816 8548
rect 5810 8508 5816 8520
rect 5868 8508 5874 8560
rect 5905 8551 5963 8557
rect 5905 8517 5917 8551
rect 5951 8548 5963 8551
rect 12710 8548 12716 8560
rect 5951 8520 12716 8548
rect 5951 8517 5963 8520
rect 5905 8511 5963 8517
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 24854 8548 24860 8560
rect 22296 8520 24860 8548
rect 22296 8489 22324 8520
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 25130 8508 25136 8560
rect 25188 8508 25194 8560
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23900 8452 23949 8480
rect 23900 8440 23906 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2832 8384 4169 8412
rect 2832 8372 2838 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 24486 8412 24492 8424
rect 23339 8384 24492 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 24486 8372 24492 8384
rect 24544 8372 24550 8424
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 16632 7840 18705 7868
rect 16632 7828 16638 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20806 7868 20812 7880
rect 20395 7840 20812 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23290 7868 23296 7880
rect 22879 7840 23296 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 20533 7803 20591 7809
rect 20533 7769 20545 7803
rect 20579 7800 20591 7803
rect 21266 7800 21272 7812
rect 20579 7772 21272 7800
rect 20579 7769 20591 7772
rect 20533 7763 20591 7769
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 23845 7803 23903 7809
rect 23845 7769 23857 7803
rect 23891 7800 23903 7803
rect 24946 7800 24952 7812
rect 23891 7772 24952 7800
rect 23891 7769 23903 7772
rect 23845 7763 23903 7769
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 18785 7735 18843 7741
rect 18785 7701 18797 7735
rect 18831 7732 18843 7735
rect 20438 7732 20444 7744
rect 18831 7704 20444 7732
rect 18831 7701 18843 7704
rect 18785 7695 18843 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 24670 7692 24676 7744
rect 24728 7692 24734 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 21269 7463 21327 7469
rect 21269 7429 21281 7463
rect 21315 7460 21327 7463
rect 25406 7460 25412 7472
rect 21315 7432 25412 7460
rect 21315 7429 21327 7432
rect 21269 7423 21327 7429
rect 25406 7420 25412 7432
rect 25464 7420 25470 7472
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20806 7392 20812 7404
rect 20303 7364 20812 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 20956 7364 22109 7392
rect 20956 7352 20962 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7392 24179 7395
rect 24578 7392 24584 7404
rect 24167 7364 24584 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22520 7296 22569 7324
rect 22520 7284 22526 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 24762 7284 24768 7336
rect 24820 7284 24826 7336
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 14550 6808 14556 6860
rect 14608 6848 14614 6860
rect 14608 6820 19656 6848
rect 14608 6808 14614 6820
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 19628 6789 19656 6820
rect 24854 6808 24860 6860
rect 24912 6808 24918 6860
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 16080 6752 18245 6780
rect 16080 6740 16086 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 20809 6783 20867 6789
rect 20809 6749 20821 6783
rect 20855 6749 20867 6783
rect 20809 6743 20867 6749
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6712 18475 6715
rect 19702 6712 19708 6724
rect 18463 6684 19708 6712
rect 18463 6681 18475 6684
rect 18417 6675 18475 6681
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 6270 6644 6276 6656
rect 3200 6616 6276 6644
rect 3200 6604 3206 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20824 6644 20852 6743
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24946 6780 24952 6792
rect 23891 6752 24952 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 23474 6672 23480 6724
rect 23532 6712 23538 6724
rect 24486 6712 24492 6724
rect 23532 6684 24492 6712
rect 23532 6672 23538 6684
rect 24486 6672 24492 6684
rect 24544 6712 24550 6724
rect 24673 6715 24731 6721
rect 24673 6712 24685 6715
rect 24544 6684 24685 6712
rect 24544 6672 24550 6684
rect 24673 6681 24685 6684
rect 24719 6681 24731 6715
rect 24673 6675 24731 6681
rect 19475 6616 20852 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 20898 6440 20904 6452
rect 19567 6412 20904 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 21269 6375 21327 6381
rect 12124 6344 20116 6372
rect 12124 6332 12130 6344
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 20088 6313 20116 6344
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 22370 6372 22376 6384
rect 21315 6344 22376 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 22370 6332 22376 6344
rect 22428 6332 22434 6384
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 17368 6276 19441 6304
rect 17368 6264 17374 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 20073 6307 20131 6313
rect 20073 6273 20085 6307
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 24118 6264 24124 6316
rect 24176 6264 24182 6316
rect 5166 6196 5172 6248
rect 5224 6236 5230 6248
rect 11238 6236 11244 6248
rect 5224 6208 11244 6236
rect 5224 6196 5230 6208
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 22186 6196 22192 6248
rect 22244 6236 22250 6248
rect 22557 6239 22615 6245
rect 22557 6236 22569 6239
rect 22244 6208 22569 6236
rect 22244 6196 22250 6208
rect 22557 6205 22569 6208
rect 22603 6205 22615 6239
rect 22557 6199 22615 6205
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 24762 6100 24768 6112
rect 20864 6072 24768 6100
rect 20864 6060 20870 6072
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 22094 5896 22100 5908
rect 20027 5868 22100 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 24762 5856 24768 5908
rect 24820 5856 24826 5908
rect 20438 5788 20444 5840
rect 20496 5828 20502 5840
rect 20496 5800 22600 5828
rect 20496 5788 20502 5800
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 21177 5763 21235 5769
rect 21177 5760 21189 5763
rect 20680 5732 21189 5760
rect 20680 5720 20686 5732
rect 21177 5729 21189 5732
rect 21223 5729 21235 5763
rect 21177 5723 21235 5729
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 8478 5692 8484 5704
rect 2096 5664 8484 5692
rect 2096 5652 2102 5664
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 22572 5701 22600 5800
rect 23017 5763 23075 5769
rect 23017 5729 23029 5763
rect 23063 5729 23075 5763
rect 23017 5723 23075 5729
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 15838 5624 15844 5636
rect 10652 5596 15844 5624
rect 10652 5584 10658 5596
rect 15838 5584 15844 5596
rect 15896 5584 15902 5636
rect 21726 5584 21732 5636
rect 21784 5624 21790 5636
rect 23032 5624 23060 5723
rect 21784 5596 23060 5624
rect 21784 5584 21790 5596
rect 24486 5584 24492 5636
rect 24544 5624 24550 5636
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 24544 5596 24685 5624
rect 24544 5584 24550 5596
rect 24673 5593 24685 5596
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 2130 5516 2136 5568
rect 2188 5556 2194 5568
rect 6454 5556 6460 5568
rect 2188 5528 6460 5556
rect 2188 5516 2194 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10318 5556 10324 5568
rect 9640 5528 10324 5556
rect 9640 5516 9646 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 23842 5556 23848 5568
rect 22796 5528 23848 5556
rect 22796 5516 22802 5528
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 18046 5216 18052 5228
rect 17911 5188 18052 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 19610 5176 19616 5228
rect 19668 5176 19674 5228
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 19760 5188 22017 5216
rect 19760 5176 19766 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5216 24179 5219
rect 24670 5216 24676 5228
rect 24167 5188 24676 5216
rect 24167 5185 24179 5188
rect 24121 5179 24179 5185
rect 24670 5176 24676 5188
rect 24728 5176 24734 5228
rect 18969 5151 19027 5157
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19426 5148 19432 5160
rect 19015 5120 19432 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19426 5108 19432 5120
rect 19484 5108 19490 5160
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19576 5120 20085 5148
rect 19576 5108 19582 5120
rect 20073 5117 20085 5120
rect 20119 5117 20131 5151
rect 20073 5111 20131 5117
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22336 5120 22477 5148
rect 22336 5108 22342 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 12618 5012 12624 5024
rect 9456 4984 12624 5012
rect 9456 4972 9462 4984
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 16117 5015 16175 5021
rect 16117 4981 16129 5015
rect 16163 5012 16175 5015
rect 23566 5012 23572 5024
rect 16163 4984 23572 5012
rect 16163 4981 16175 4984
rect 16117 4975 16175 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 6362 4808 6368 4820
rect 3292 4780 6368 4808
rect 3292 4768 3298 4780
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 11606 4808 11612 4820
rect 6512 4780 11612 4808
rect 6512 4768 6518 4780
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 25314 4768 25320 4820
rect 25372 4768 25378 4820
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 23477 4675 23535 4681
rect 23477 4672 23489 4675
rect 18104 4644 23489 4672
rect 18104 4632 18110 4644
rect 23477 4641 23489 4644
rect 23523 4641 23535 4675
rect 23477 4635 23535 4641
rect 17494 4564 17500 4616
rect 17552 4564 17558 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 20530 4564 20536 4616
rect 20588 4604 20594 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 20588 4576 21281 4604
rect 20588 4564 20594 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 23201 4607 23259 4613
rect 23201 4604 23213 4607
rect 21269 4567 21327 4573
rect 22664 4576 23213 4604
rect 18322 4496 18328 4548
rect 18380 4496 18386 4548
rect 20346 4496 20352 4548
rect 20404 4496 20410 4548
rect 21082 4496 21088 4548
rect 21140 4536 21146 4548
rect 22189 4539 22247 4545
rect 22189 4536 22201 4539
rect 21140 4508 22201 4536
rect 21140 4496 21146 4508
rect 22189 4505 22201 4508
rect 22235 4505 22247 4539
rect 22189 4499 22247 4505
rect 19794 4428 19800 4480
rect 19852 4468 19858 4480
rect 22664 4468 22692 4576
rect 23201 4573 23213 4576
rect 23247 4604 23259 4607
rect 23750 4604 23756 4616
rect 23247 4576 23756 4604
rect 23247 4573 23259 4576
rect 23201 4567 23259 4573
rect 23750 4564 23756 4576
rect 23808 4564 23814 4616
rect 19852 4440 22692 4468
rect 19852 4428 19858 4440
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 8938 4196 8944 4208
rect 5132 4168 8944 4196
rect 5132 4156 5138 4168
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 11514 4156 11520 4208
rect 11572 4196 11578 4208
rect 13722 4196 13728 4208
rect 11572 4168 13728 4196
rect 11572 4156 11578 4168
rect 13722 4156 13728 4168
rect 13780 4156 13786 4208
rect 21542 4156 21548 4208
rect 21600 4196 21606 4208
rect 21600 4168 22140 4196
rect 21600 4156 21606 4168
rect 1118 4088 1124 4140
rect 1176 4128 1182 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1176 4100 1777 4128
rect 1176 4088 1182 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4128 7895 4131
rect 8846 4128 8852 4140
rect 7883 4100 8852 4128
rect 7883 4097 7895 4100
rect 7837 4091 7895 4097
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13630 4128 13636 4140
rect 13219 4100 13636 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13630 4088 13636 4100
rect 13688 4088 13694 4140
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 15252 4100 16865 4128
rect 15252 4088 15258 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 22112 4137 22140 4168
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 12860 4032 13461 4060
rect 12860 4020 12866 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18472 4032 19165 4060
rect 18472 4020 18478 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20312 4032 22477 4060
rect 20312 4020 20318 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 5534 3992 5540 4004
rect 1627 3964 5540 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 7834 3952 7840 4004
rect 7892 3992 7898 4004
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7892 3964 8033 3992
rect 7892 3952 7898 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 9490 3952 9496 4004
rect 9548 3952 9554 4004
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 24320 3992 24348 4023
rect 21600 3964 24348 3992
rect 21600 3952 21606 3964
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2774 3720 2780 3732
rect 2363 3692 2780 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3418 3720 3424 3732
rect 3283 3692 3424 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5074 3680 5080 3732
rect 5132 3680 5138 3732
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6730 3720 6736 3732
rect 6595 3692 6736 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7650 3680 7656 3732
rect 7708 3680 7714 3732
rect 8386 3680 8392 3732
rect 8444 3680 8450 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 11514 3680 11520 3732
rect 11572 3680 11578 3732
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 4982 3652 4988 3664
rect 1903 3624 4988 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 5629 3655 5687 3661
rect 5629 3621 5641 3655
rect 5675 3652 5687 3655
rect 16022 3652 16028 3664
rect 5675 3624 16028 3652
rect 5675 3621 5687 3624
rect 5629 3615 5687 3621
rect 16022 3612 16028 3624
rect 16080 3612 16086 3664
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12584 3556 12817 3584
rect 12584 3544 12590 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17736 3556 19901 3584
rect 17736 3544 17742 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21358 3544 21364 3596
rect 21416 3584 21422 3596
rect 23290 3584 23296 3596
rect 21416 3556 23296 3584
rect 21416 3544 21422 3556
rect 23290 3544 23296 3556
rect 23348 3544 23354 3596
rect 23474 3544 23480 3596
rect 23532 3544 23538 3596
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2774 3516 2780 3528
rect 2547 3488 2780 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2924 3488 3065 3516
rect 2924 3476 2930 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4856 3488 4905 3516
rect 4856 3476 4862 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5592 3488 5825 3516
rect 5592 3476 5598 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 5813 3479 5871 3485
rect 6270 3476 6276 3528
rect 6328 3516 6334 3528
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 6328 3488 6377 3516
rect 6328 3476 6334 3488
rect 6365 3485 6377 3488
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7469 3519 7527 3525
rect 7469 3516 7481 3519
rect 7432 3488 7481 3516
rect 7432 3476 7438 3488
rect 7469 3485 7481 3488
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7892 3488 8217 3516
rect 7892 3476 7898 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9582 3516 9588 3528
rect 9355 3488 9588 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 10008 3488 10057 3516
rect 10008 3476 10014 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 1544 3420 1685 3448
rect 1544 3408 1550 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 1673 3411 1731 3417
rect 10336 3380 10364 3479
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 10744 3488 11345 3516
rect 10744 3476 10750 3488
rect 11333 3485 11345 3488
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12452 3448 12480 3479
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 16114 3476 16120 3528
rect 16172 3476 16178 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17828 3488 19441 3516
rect 17828 3476 17834 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21266 3476 21272 3528
rect 21324 3476 21330 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 14458 3448 14464 3460
rect 12452 3420 14464 3448
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 22189 3451 22247 3457
rect 22189 3448 22201 3451
rect 19208 3420 22201 3448
rect 19208 3408 19214 3420
rect 22189 3417 22201 3420
rect 22235 3417 22247 3451
rect 23216 3448 23244 3479
rect 24302 3448 24308 3460
rect 23216 3420 24308 3448
rect 22189 3411 22247 3417
rect 24302 3408 24308 3420
rect 24360 3408 24366 3460
rect 14734 3380 14740 3392
rect 10336 3352 14740 3380
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22830 3380 22836 3392
rect 22060 3352 22836 3380
rect 22060 3340 22066 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2130 3136 2136 3188
rect 2188 3136 2194 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 23750 3136 23756 3188
rect 23808 3176 23814 3188
rect 24857 3179 24915 3185
rect 24857 3176 24869 3179
rect 23808 3148 24869 3176
rect 23808 3136 23814 3148
rect 24857 3145 24869 3148
rect 24903 3145 24915 3179
rect 24857 3139 24915 3145
rect 3053 3111 3111 3117
rect 3053 3077 3065 3111
rect 3099 3108 3111 3111
rect 3878 3108 3884 3120
rect 3099 3080 3884 3108
rect 3099 3077 3111 3080
rect 3053 3071 3111 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3108 6055 3111
rect 6086 3108 6092 3120
rect 6043 3080 6092 3108
rect 6043 3077 6055 3080
rect 5997 3071 6055 3077
rect 6086 3068 6092 3080
rect 6144 3068 6150 3120
rect 15010 3108 15016 3120
rect 7392 3080 15016 3108
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1912 3012 1961 3040
rect 1912 3000 1918 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3326 3040 3332 3052
rect 2915 3012 3332 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3694 3040 3700 3052
rect 3559 3012 3700 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4430 3040 4436 3052
rect 4295 3012 4436 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5166 3040 5172 3052
rect 5031 3012 5172 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5902 3040 5908 3052
rect 5859 3012 5908 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 7392 3049 7420 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 23934 3108 23940 3120
rect 19484 3080 23940 3108
rect 19484 3068 19490 3080
rect 23934 3068 23940 3080
rect 23992 3068 23998 3120
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 9398 3040 9404 3052
rect 8895 3012 9404 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 10594 3000 10600 3052
rect 10652 3000 10658 3052
rect 11974 3000 11980 3052
rect 12032 3000 12038 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12492 3012 13001 3040
rect 12492 3000 12498 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 16666 3000 16672 3052
rect 16724 3040 16730 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16724 3012 16865 3040
rect 16724 3000 16730 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18693 3043 18751 3049
rect 18693 3040 18705 3043
rect 17920 3012 18705 3040
rect 17920 3000 17926 3012
rect 18693 3009 18705 3012
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 7064 2944 7113 2972
rect 7064 2932 7070 2944
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 7101 2935 7159 2941
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 8536 2944 8585 2972
rect 8536 2932 8542 2944
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8573 2935 8631 2941
rect 10318 2932 10324 2984
rect 10376 2932 10382 2984
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 11790 2972 11796 2984
rect 11747 2944 11796 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2972 22615 2975
rect 24486 2972 24492 2984
rect 22603 2944 24492 2972
rect 22603 2941 22615 2944
rect 22557 2935 22615 2941
rect 3697 2907 3755 2913
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 7282 2904 7288 2916
rect 3743 2876 7288 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 19168 2904 19196 2935
rect 16632 2876 19196 2904
rect 16632 2864 16638 2876
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 21082 2904 21088 2916
rect 19944 2876 21088 2904
rect 19944 2864 19950 2876
rect 21082 2864 21088 2876
rect 21140 2864 21146 2916
rect 22296 2904 22324 2935
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 25038 2904 25044 2916
rect 22296 2876 25044 2904
rect 25038 2864 25044 2876
rect 25096 2864 25102 2916
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 5074 2836 5080 2848
rect 4479 2808 5080 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 11054 2836 11060 2848
rect 9548 2808 11060 2836
rect 9548 2796 9554 2808
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 18322 2836 18328 2848
rect 17368 2808 18328 2836
rect 17368 2796 17374 2808
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 20346 2836 20352 2848
rect 18840 2808 20352 2836
rect 18840 2796 18846 2808
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 22278 2836 22284 2848
rect 21048 2808 22284 2836
rect 21048 2796 21054 2808
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 2038 2592 2044 2644
rect 2096 2592 2102 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6454 2632 6460 2644
rect 5951 2604 6460 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 10778 2632 10784 2644
rect 6886 2604 10784 2632
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 6886 2496 6914 2604
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 15286 2632 15292 2644
rect 11747 2604 15292 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 8662 2564 8668 2576
rect 7331 2536 8668 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 15930 2564 15936 2576
rect 9692 2536 15936 2564
rect 4479 2468 6914 2496
rect 7745 2499 7803 2505
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 9490 2496 9496 2508
rect 7791 2468 9496 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2222 2428 2228 2440
rect 1903 2400 2228 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2648 2400 2789 2428
rect 2648 2388 2654 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 2777 2391 2835 2397
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 4120 2400 4169 2428
rect 4120 2388 4126 2400
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6638 2428 6644 2440
rect 5767 2400 6644 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 8021 2431 8079 2437
rect 6886 2400 7880 2428
rect 6886 2360 6914 2400
rect 2608 2332 6914 2360
rect 7101 2363 7159 2369
rect 2608 2301 2636 2332
rect 7101 2329 7113 2363
rect 7147 2360 7159 2363
rect 7852 2360 7880 2400
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 9692 2428 9720 2536
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11756 2468 12388 2496
rect 11756 2456 11762 2468
rect 8067 2400 9720 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 12360 2437 12388 2468
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15160 2468 17325 2496
rect 15160 2456 15166 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 17313 2459 17371 2465
rect 18156 2468 19901 2496
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11480 2400 11897 2428
rect 11480 2388 11486 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 16298 2428 16304 2440
rect 14691 2400 16304 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 18156 2428 18184 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 17000 2400 18184 2428
rect 18248 2400 19441 2428
rect 17000 2388 17006 2400
rect 9030 2360 9036 2372
rect 7147 2332 7788 2360
rect 7852 2332 9036 2360
rect 7147 2329 7159 2332
rect 7101 2323 7159 2329
rect 7760 2304 7788 2332
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 10965 2363 11023 2369
rect 10965 2329 10977 2363
rect 11011 2360 11023 2363
rect 12158 2360 12164 2372
rect 11011 2332 12164 2360
rect 11011 2329 11023 2332
rect 10965 2323 11023 2329
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 17034 2320 17040 2372
rect 17092 2360 17098 2372
rect 18248 2360 18276 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21508 2400 22017 2428
rect 21508 2388 21514 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 17092 2332 18276 2360
rect 17092 2320 17098 2332
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 22480 2360 22508 2459
rect 18564 2332 22508 2360
rect 18564 2320 18570 2332
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2261 2651 2295
rect 2593 2255 2651 2261
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 5356 54204 5408 54256
rect 6828 54204 6880 54256
rect 9404 54204 9456 54256
rect 10876 54247 10928 54256
rect 10876 54213 10885 54247
rect 10885 54213 10919 54247
rect 10919 54213 10928 54247
rect 10876 54204 10928 54213
rect 14924 54204 14976 54256
rect 16028 54204 16080 54256
rect 4712 54136 4764 54188
rect 7472 54136 7524 54188
rect 9864 54179 9916 54188
rect 9864 54145 9873 54179
rect 9873 54145 9907 54179
rect 9907 54145 9916 54179
rect 9864 54136 9916 54145
rect 12072 54179 12124 54188
rect 12072 54145 12081 54179
rect 12081 54145 12115 54179
rect 12115 54145 12124 54179
rect 12072 54136 12124 54145
rect 14556 54136 14608 54188
rect 15292 54136 15344 54188
rect 17132 54204 17184 54256
rect 19340 54204 19392 54256
rect 17500 54136 17552 54188
rect 18604 54136 18656 54188
rect 20076 54204 20128 54256
rect 24124 54204 24176 54256
rect 21180 54136 21232 54188
rect 8576 54068 8628 54120
rect 11980 54068 12032 54120
rect 22744 54136 22796 54188
rect 23756 54068 23808 54120
rect 15752 54000 15804 54052
rect 20628 54000 20680 54052
rect 14832 53975 14884 53984
rect 14832 53941 14841 53975
rect 14841 53941 14875 53975
rect 14875 53941 14884 53975
rect 14832 53932 14884 53941
rect 15568 53975 15620 53984
rect 15568 53941 15577 53975
rect 15577 53941 15611 53975
rect 15611 53941 15620 53975
rect 15568 53932 15620 53941
rect 16120 53975 16172 53984
rect 16120 53941 16129 53975
rect 16129 53941 16163 53975
rect 16163 53941 16172 53975
rect 16120 53932 16172 53941
rect 17776 53975 17828 53984
rect 17776 53941 17785 53975
rect 17785 53941 17819 53975
rect 17819 53941 17828 53975
rect 17776 53932 17828 53941
rect 18512 53975 18564 53984
rect 18512 53941 18521 53975
rect 18521 53941 18555 53975
rect 18555 53941 18564 53975
rect 18512 53932 18564 53941
rect 19616 53975 19668 53984
rect 19616 53941 19625 53975
rect 19625 53941 19659 53975
rect 19659 53941 19668 53975
rect 19616 53932 19668 53941
rect 20996 53932 21048 53984
rect 21824 53932 21876 53984
rect 23388 53932 23440 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 4620 53592 4672 53644
rect 7564 53592 7616 53644
rect 8300 53635 8352 53644
rect 8300 53601 8309 53635
rect 8309 53601 8343 53635
rect 8343 53601 8352 53635
rect 8300 53592 8352 53601
rect 9036 53592 9088 53644
rect 9680 53592 9732 53644
rect 10508 53635 10560 53644
rect 10508 53601 10517 53635
rect 10517 53601 10551 53635
rect 10551 53601 10560 53635
rect 10508 53592 10560 53601
rect 11612 53592 11664 53644
rect 25596 53592 25648 53644
rect 5448 53567 5500 53576
rect 5448 53533 5457 53567
rect 5457 53533 5491 53567
rect 5491 53533 5500 53567
rect 5448 53524 5500 53533
rect 7380 53567 7432 53576
rect 7380 53533 7389 53567
rect 7389 53533 7423 53567
rect 7423 53533 7432 53567
rect 7380 53524 7432 53533
rect 10048 53567 10100 53576
rect 10048 53533 10057 53567
rect 10057 53533 10091 53567
rect 10091 53533 10100 53567
rect 10048 53524 10100 53533
rect 11704 53567 11756 53576
rect 11704 53533 11713 53567
rect 11713 53533 11747 53567
rect 11747 53533 11756 53567
rect 11704 53524 11756 53533
rect 13820 53524 13872 53576
rect 14188 53524 14240 53576
rect 15660 53524 15712 53576
rect 16396 53524 16448 53576
rect 16764 53524 16816 53576
rect 17868 53524 17920 53576
rect 18328 53524 18380 53576
rect 18972 53524 19024 53576
rect 20444 53524 20496 53576
rect 20812 53524 20864 53576
rect 21548 53524 21600 53576
rect 6644 53456 6696 53508
rect 18420 53456 18472 53508
rect 23296 53524 23348 53576
rect 12532 53388 12584 53440
rect 14464 53431 14516 53440
rect 14464 53397 14473 53431
rect 14473 53397 14507 53431
rect 14507 53397 14516 53431
rect 14464 53388 14516 53397
rect 15936 53431 15988 53440
rect 15936 53397 15945 53431
rect 15945 53397 15979 53431
rect 15979 53397 15988 53431
rect 15936 53388 15988 53397
rect 16212 53388 16264 53440
rect 17224 53431 17276 53440
rect 17224 53397 17233 53431
rect 17233 53397 17267 53431
rect 17267 53397 17276 53431
rect 17224 53388 17276 53397
rect 18696 53431 18748 53440
rect 18696 53397 18705 53431
rect 18705 53397 18739 53431
rect 18739 53397 18748 53431
rect 18696 53388 18748 53397
rect 20076 53388 20128 53440
rect 25872 53456 25924 53508
rect 21456 53431 21508 53440
rect 21456 53397 21465 53431
rect 21465 53397 21499 53431
rect 21499 53397 21508 53431
rect 21456 53388 21508 53397
rect 21548 53388 21600 53440
rect 22008 53431 22060 53440
rect 22008 53397 22017 53431
rect 22017 53397 22051 53431
rect 22051 53397 22060 53431
rect 22008 53388 22060 53397
rect 23296 53388 23348 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 2780 53184 2832 53236
rect 4252 53116 4304 53168
rect 5724 53159 5776 53168
rect 5724 53125 5733 53159
rect 5733 53125 5767 53159
rect 5767 53125 5776 53159
rect 5724 53116 5776 53125
rect 12716 53116 12768 53168
rect 24860 53159 24912 53168
rect 24860 53125 24869 53159
rect 24869 53125 24903 53159
rect 24903 53125 24912 53159
rect 24860 53116 24912 53125
rect 6368 53048 6420 53100
rect 6828 53091 6880 53100
rect 6828 53057 6837 53091
rect 6837 53057 6871 53091
rect 6871 53057 6880 53091
rect 6828 53048 6880 53057
rect 9220 53048 9272 53100
rect 9404 53048 9456 53100
rect 10508 53048 10560 53100
rect 13452 53048 13504 53100
rect 19708 53048 19760 53100
rect 21916 53048 21968 53100
rect 22284 53048 22336 53100
rect 25964 53048 26016 53100
rect 6552 52980 6604 53032
rect 8668 53023 8720 53032
rect 8668 52989 8677 53023
rect 8677 52989 8711 53023
rect 8711 52989 8720 53023
rect 8668 52980 8720 52989
rect 10140 52980 10192 53032
rect 11244 52980 11296 53032
rect 14556 52955 14608 52964
rect 14556 52921 14565 52955
rect 14565 52921 14599 52955
rect 14599 52921 14608 52955
rect 14556 52912 14608 52921
rect 3976 52844 4028 52896
rect 4252 52844 4304 52896
rect 13728 52887 13780 52896
rect 13728 52853 13737 52887
rect 13737 52853 13771 52887
rect 13771 52853 13780 52887
rect 13728 52844 13780 52853
rect 19800 52887 19852 52896
rect 19800 52853 19809 52887
rect 19809 52853 19843 52887
rect 19843 52853 19852 52887
rect 19800 52844 19852 52853
rect 22192 52887 22244 52896
rect 22192 52853 22201 52887
rect 22201 52853 22235 52887
rect 22235 52853 22244 52887
rect 22192 52844 22244 52853
rect 22744 52887 22796 52896
rect 22744 52853 22753 52887
rect 22753 52853 22787 52887
rect 22787 52853 22796 52887
rect 22744 52844 22796 52853
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 2044 52640 2096 52692
rect 3424 52640 3476 52692
rect 12072 52640 12124 52692
rect 23756 52683 23808 52692
rect 23756 52649 23765 52683
rect 23765 52649 23799 52683
rect 23799 52649 23808 52683
rect 23756 52640 23808 52649
rect 940 52572 992 52624
rect 4436 52572 4488 52624
rect 13452 52572 13504 52624
rect 1308 52504 1360 52556
rect 6000 52504 6052 52556
rect 6092 52547 6144 52556
rect 6092 52513 6101 52547
rect 6101 52513 6135 52547
rect 6135 52513 6144 52547
rect 6092 52504 6144 52513
rect 7840 52547 7892 52556
rect 7840 52513 7849 52547
rect 7849 52513 7883 52547
rect 7883 52513 7892 52547
rect 7840 52504 7892 52513
rect 9772 52504 9824 52556
rect 3148 52436 3200 52488
rect 3332 52436 3384 52488
rect 5724 52436 5776 52488
rect 6460 52436 6512 52488
rect 6920 52436 6972 52488
rect 8944 52436 8996 52488
rect 9588 52436 9640 52488
rect 11980 52479 12032 52488
rect 11980 52445 11989 52479
rect 11989 52445 12023 52479
rect 12023 52445 12032 52479
rect 11980 52436 12032 52445
rect 12348 52436 12400 52488
rect 13360 52436 13412 52488
rect 14096 52436 14148 52488
rect 24492 52436 24544 52488
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 11704 52139 11756 52148
rect 11704 52105 11713 52139
rect 11713 52105 11747 52139
rect 11747 52105 11756 52139
rect 11704 52096 11756 52105
rect 5632 52028 5684 52080
rect 6276 51960 6328 52012
rect 7104 52003 7156 52012
rect 7104 51969 7113 52003
rect 7113 51969 7147 52003
rect 7147 51969 7156 52003
rect 7104 51960 7156 51969
rect 9128 52003 9180 52012
rect 9128 51969 9137 52003
rect 9137 51969 9171 52003
rect 9171 51969 9180 52003
rect 9128 51960 9180 51969
rect 11888 52003 11940 52012
rect 11888 51969 11897 52003
rect 11897 51969 11931 52003
rect 11931 51969 11940 52003
rect 11888 51960 11940 51969
rect 25136 52003 25188 52012
rect 25136 51969 25145 52003
rect 25145 51969 25179 52003
rect 25179 51969 25188 52003
rect 25136 51960 25188 51969
rect 3516 51935 3568 51944
rect 3516 51901 3525 51935
rect 3525 51901 3559 51935
rect 3559 51901 3568 51935
rect 3516 51892 3568 51901
rect 4988 51892 5040 51944
rect 7012 51892 7064 51944
rect 9680 51935 9732 51944
rect 9680 51901 9689 51935
rect 9689 51901 9723 51935
rect 9723 51901 9732 51935
rect 9680 51892 9732 51901
rect 24124 51756 24176 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 4712 51552 4764 51604
rect 2780 51459 2832 51468
rect 2780 51425 2789 51459
rect 2789 51425 2823 51459
rect 2823 51425 2832 51459
rect 2780 51416 2832 51425
rect 4160 51416 4212 51468
rect 6920 51416 6972 51468
rect 4252 51348 4304 51400
rect 7288 51348 7340 51400
rect 25044 51391 25096 51400
rect 25044 51357 25053 51391
rect 25053 51357 25087 51391
rect 25087 51357 25096 51391
rect 25044 51348 25096 51357
rect 7012 51280 7064 51332
rect 5540 51212 5592 51264
rect 25596 51212 25648 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 5540 51008 5592 51060
rect 9864 51051 9916 51060
rect 9864 51017 9873 51051
rect 9873 51017 9907 51051
rect 9907 51017 9916 51051
rect 9864 51008 9916 51017
rect 10508 51051 10560 51060
rect 10508 51017 10517 51051
rect 10517 51017 10551 51051
rect 10551 51017 10560 51051
rect 10508 51008 10560 51017
rect 3700 50872 3752 50924
rect 7196 50872 7248 50924
rect 8392 50872 8444 50924
rect 9956 50872 10008 50924
rect 25044 50915 25096 50924
rect 25044 50881 25053 50915
rect 25053 50881 25087 50915
rect 25087 50881 25096 50915
rect 25044 50872 25096 50881
rect 940 50804 992 50856
rect 2872 50804 2924 50856
rect 7564 50736 7616 50788
rect 25688 50668 25740 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 7104 50464 7156 50516
rect 9404 50439 9456 50448
rect 9404 50405 9413 50439
rect 9413 50405 9447 50439
rect 9447 50405 9456 50439
rect 9404 50396 9456 50405
rect 3424 50328 3476 50380
rect 4436 50371 4488 50380
rect 4436 50337 4445 50371
rect 4445 50337 4479 50371
rect 4479 50337 4488 50371
rect 4436 50328 4488 50337
rect 3516 50260 3568 50312
rect 5540 50260 5592 50312
rect 6920 50260 6972 50312
rect 25044 50303 25096 50312
rect 25044 50269 25053 50303
rect 25053 50269 25087 50303
rect 25087 50269 25096 50303
rect 25044 50260 25096 50269
rect 10416 50192 10468 50244
rect 25780 50124 25832 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 7380 49920 7432 49972
rect 9588 49895 9640 49904
rect 9588 49861 9597 49895
rect 9597 49861 9631 49895
rect 9631 49861 9640 49895
rect 9588 49852 9640 49861
rect 1768 49827 1820 49836
rect 1768 49793 1777 49827
rect 1777 49793 1811 49827
rect 1811 49793 1820 49827
rect 1768 49784 1820 49793
rect 7104 49784 7156 49836
rect 9312 49784 9364 49836
rect 1676 49716 1728 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 1216 49240 1268 49292
rect 1584 49215 1636 49224
rect 1584 49181 1593 49215
rect 1593 49181 1627 49215
rect 1627 49181 1636 49215
rect 1584 49172 1636 49181
rect 25044 49215 25096 49224
rect 25044 49181 25053 49215
rect 25053 49181 25087 49215
rect 25087 49181 25096 49215
rect 25044 49172 25096 49181
rect 21456 49036 21508 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 11980 48832 12032 48884
rect 3976 48764 4028 48816
rect 11704 48696 11756 48748
rect 25044 48739 25096 48748
rect 25044 48705 25053 48739
rect 25053 48705 25087 48739
rect 25087 48705 25096 48739
rect 25044 48696 25096 48705
rect 9772 48628 9824 48680
rect 10784 48560 10836 48612
rect 9404 48492 9456 48544
rect 25136 48492 25188 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 25044 48127 25096 48136
rect 25044 48093 25053 48127
rect 25053 48093 25087 48127
rect 25087 48093 25096 48127
rect 25044 48084 25096 48093
rect 940 48016 992 48068
rect 3884 48016 3936 48068
rect 25412 47948 25464 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 25044 47651 25096 47660
rect 25044 47617 25053 47651
rect 25053 47617 25087 47651
rect 25087 47617 25096 47651
rect 25044 47608 25096 47617
rect 21364 47404 21416 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 6828 47200 6880 47252
rect 11888 47200 11940 47252
rect 17408 47200 17460 47252
rect 16396 47132 16448 47184
rect 15752 47064 15804 47116
rect 16120 47064 16172 47116
rect 10600 46996 10652 47048
rect 11612 46996 11664 47048
rect 15016 46860 15068 46912
rect 16764 46928 16816 46980
rect 16948 46928 17000 46980
rect 17776 46971 17828 46980
rect 17776 46937 17785 46971
rect 17785 46937 17819 46971
rect 17819 46937 17828 46971
rect 17776 46928 17828 46937
rect 17316 46903 17368 46912
rect 17316 46869 17325 46903
rect 17325 46869 17359 46903
rect 17359 46869 17368 46903
rect 17316 46860 17368 46869
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7012 46699 7064 46708
rect 7012 46665 7021 46699
rect 7021 46665 7055 46699
rect 7055 46665 7064 46699
rect 7012 46656 7064 46665
rect 15384 46699 15436 46708
rect 15384 46665 15393 46699
rect 15393 46665 15427 46699
rect 15427 46665 15436 46699
rect 15384 46656 15436 46665
rect 16396 46656 16448 46708
rect 17224 46699 17276 46708
rect 17224 46665 17233 46699
rect 17233 46665 17267 46699
rect 17267 46665 17276 46699
rect 17224 46656 17276 46665
rect 18696 46656 18748 46708
rect 18880 46588 18932 46640
rect 7840 46520 7892 46572
rect 15016 46520 15068 46572
rect 18420 46563 18472 46572
rect 18420 46529 18429 46563
rect 18429 46529 18463 46563
rect 18463 46529 18472 46563
rect 18420 46520 18472 46529
rect 18512 46520 18564 46572
rect 13360 46452 13412 46504
rect 16028 46452 16080 46504
rect 17408 46495 17460 46504
rect 17408 46461 17417 46495
rect 17417 46461 17451 46495
rect 17451 46461 17460 46495
rect 17408 46452 17460 46461
rect 18696 46495 18748 46504
rect 18696 46461 18705 46495
rect 18705 46461 18739 46495
rect 18739 46461 18748 46495
rect 18696 46452 18748 46461
rect 17224 46316 17276 46368
rect 17868 46316 17920 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 5724 46112 5776 46164
rect 17408 46112 17460 46164
rect 22468 46044 22520 46096
rect 17592 45976 17644 46028
rect 19800 45976 19852 46028
rect 19984 46019 20036 46028
rect 19984 45985 19993 46019
rect 19993 45985 20027 46019
rect 20027 45985 20036 46019
rect 19984 45976 20036 45985
rect 22100 45976 22152 46028
rect 940 45908 992 45960
rect 9680 45908 9732 45960
rect 9864 45908 9916 45960
rect 15844 45951 15896 45960
rect 15844 45917 15853 45951
rect 15853 45917 15887 45951
rect 15887 45917 15896 45951
rect 15844 45908 15896 45917
rect 22008 45908 22060 45960
rect 24676 45908 24728 45960
rect 7288 45840 7340 45892
rect 16580 45840 16632 45892
rect 19616 45772 19668 45824
rect 19800 45815 19852 45824
rect 19800 45781 19809 45815
rect 19809 45781 19843 45815
rect 19843 45781 19852 45815
rect 19800 45772 19852 45781
rect 20628 45772 20680 45824
rect 22376 45772 22428 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 7196 45500 7248 45552
rect 15844 45568 15896 45620
rect 7656 45432 7708 45484
rect 10232 45432 10284 45484
rect 13636 45500 13688 45552
rect 15016 45500 15068 45552
rect 18512 45500 18564 45552
rect 19156 45500 19208 45552
rect 20076 45543 20128 45552
rect 20076 45509 20085 45543
rect 20085 45509 20119 45543
rect 20119 45509 20128 45543
rect 20076 45500 20128 45509
rect 21824 45500 21876 45552
rect 11796 45475 11848 45484
rect 11796 45441 11805 45475
rect 11805 45441 11839 45475
rect 11839 45441 11848 45475
rect 11796 45432 11848 45441
rect 16856 45475 16908 45484
rect 16856 45441 16865 45475
rect 16865 45441 16899 45475
rect 16899 45441 16908 45475
rect 16856 45432 16908 45441
rect 24584 45432 24636 45484
rect 7472 45364 7524 45416
rect 13360 45407 13412 45416
rect 13360 45373 13369 45407
rect 13369 45373 13403 45407
rect 13403 45373 13412 45407
rect 13360 45364 13412 45373
rect 15384 45364 15436 45416
rect 18696 45364 18748 45416
rect 20352 45407 20404 45416
rect 20352 45373 20361 45407
rect 20361 45373 20395 45407
rect 20395 45373 20404 45407
rect 20352 45364 20404 45373
rect 24768 45407 24820 45416
rect 24768 45373 24777 45407
rect 24777 45373 24811 45407
rect 24811 45373 24820 45407
rect 24768 45364 24820 45373
rect 8392 45339 8444 45348
rect 8392 45305 8401 45339
rect 8401 45305 8435 45339
rect 8435 45305 8444 45339
rect 8392 45296 8444 45305
rect 9956 45296 10008 45348
rect 15108 45271 15160 45280
rect 15108 45237 15117 45271
rect 15117 45237 15151 45271
rect 15151 45237 15160 45271
rect 15108 45228 15160 45237
rect 18604 45271 18656 45280
rect 18604 45237 18613 45271
rect 18613 45237 18647 45271
rect 18647 45237 18656 45271
rect 18604 45228 18656 45237
rect 19708 45271 19760 45280
rect 19708 45237 19717 45271
rect 19717 45237 19751 45271
rect 19751 45237 19760 45271
rect 19708 45228 19760 45237
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 6368 45024 6420 45076
rect 9128 45024 9180 45076
rect 16028 45067 16080 45076
rect 16028 45033 16037 45067
rect 16037 45033 16071 45067
rect 16071 45033 16080 45067
rect 16028 45024 16080 45033
rect 16396 45024 16448 45076
rect 24584 45067 24636 45076
rect 24584 45033 24593 45067
rect 24593 45033 24627 45067
rect 24627 45033 24636 45067
rect 24584 45024 24636 45033
rect 21916 44888 21968 44940
rect 23296 44931 23348 44940
rect 23296 44897 23305 44931
rect 23305 44897 23339 44931
rect 23339 44897 23348 44931
rect 23296 44888 23348 44897
rect 23480 44931 23532 44940
rect 23480 44897 23489 44931
rect 23489 44897 23523 44931
rect 23523 44897 23532 44931
rect 23480 44888 23532 44897
rect 10692 44863 10744 44872
rect 10692 44829 10701 44863
rect 10701 44829 10735 44863
rect 10735 44829 10744 44863
rect 10692 44820 10744 44829
rect 14280 44863 14332 44872
rect 14280 44829 14289 44863
rect 14289 44829 14323 44863
rect 14323 44829 14332 44863
rect 14280 44820 14332 44829
rect 19432 44863 19484 44872
rect 19432 44829 19441 44863
rect 19441 44829 19475 44863
rect 19475 44829 19484 44863
rect 19432 44820 19484 44829
rect 21272 44820 21324 44872
rect 23848 44820 23900 44872
rect 24492 44820 24544 44872
rect 7564 44752 7616 44804
rect 10876 44752 10928 44804
rect 11060 44752 11112 44804
rect 9956 44684 10008 44736
rect 10784 44684 10836 44736
rect 14556 44795 14608 44804
rect 14556 44761 14565 44795
rect 14565 44761 14599 44795
rect 14599 44761 14608 44795
rect 14556 44752 14608 44761
rect 12348 44684 12400 44736
rect 13820 44684 13872 44736
rect 15016 44752 15068 44804
rect 19800 44752 19852 44804
rect 19984 44752 20036 44804
rect 20996 44752 21048 44804
rect 21548 44752 21600 44804
rect 23388 44752 23440 44804
rect 19340 44684 19392 44736
rect 21640 44727 21692 44736
rect 21640 44693 21649 44727
rect 21649 44693 21683 44727
rect 21683 44693 21692 44727
rect 21640 44684 21692 44693
rect 22836 44727 22888 44736
rect 22836 44693 22845 44727
rect 22845 44693 22879 44727
rect 22879 44693 22888 44727
rect 22836 44684 22888 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 6276 44480 6328 44532
rect 8668 44523 8720 44532
rect 8668 44489 8677 44523
rect 8677 44489 8711 44523
rect 8711 44489 8720 44523
rect 8668 44480 8720 44489
rect 11704 44523 11756 44532
rect 11704 44489 11713 44523
rect 11713 44489 11747 44523
rect 11747 44489 11756 44523
rect 11704 44480 11756 44489
rect 12532 44480 12584 44532
rect 15476 44480 15528 44532
rect 16212 44480 16264 44532
rect 18696 44480 18748 44532
rect 20904 44480 20956 44532
rect 21548 44480 21600 44532
rect 9956 44412 10008 44464
rect 18512 44412 18564 44464
rect 7196 44387 7248 44396
rect 7196 44353 7205 44387
rect 7205 44353 7239 44387
rect 7239 44353 7248 44387
rect 7196 44344 7248 44353
rect 7748 44344 7800 44396
rect 9036 44344 9088 44396
rect 9404 44387 9456 44396
rect 9404 44353 9413 44387
rect 9413 44353 9447 44387
rect 9447 44353 9456 44387
rect 9404 44344 9456 44353
rect 11980 44344 12032 44396
rect 12716 44344 12768 44396
rect 16856 44344 16908 44396
rect 9772 44276 9824 44328
rect 10048 44276 10100 44328
rect 10140 44276 10192 44328
rect 6920 44208 6972 44260
rect 12164 44319 12216 44328
rect 12164 44285 12173 44319
rect 12173 44285 12207 44319
rect 12207 44285 12216 44319
rect 12164 44276 12216 44285
rect 12348 44319 12400 44328
rect 12348 44285 12357 44319
rect 12357 44285 12391 44319
rect 12391 44285 12400 44319
rect 12348 44276 12400 44285
rect 14924 44276 14976 44328
rect 19524 44276 19576 44328
rect 9772 44140 9824 44192
rect 10232 44140 10284 44192
rect 11060 44140 11112 44192
rect 12256 44140 12308 44192
rect 14188 44183 14240 44192
rect 14188 44149 14197 44183
rect 14197 44149 14231 44183
rect 14231 44149 14240 44183
rect 14188 44140 14240 44149
rect 14556 44140 14608 44192
rect 16764 44140 16816 44192
rect 17408 44140 17460 44192
rect 18420 44140 18472 44192
rect 23848 44412 23900 44464
rect 24860 44344 24912 44396
rect 25320 44387 25372 44396
rect 25320 44353 25329 44387
rect 25329 44353 25363 44387
rect 25363 44353 25372 44387
rect 25320 44344 25372 44353
rect 22008 44319 22060 44328
rect 22008 44285 22017 44319
rect 22017 44285 22051 44319
rect 22051 44285 22060 44319
rect 22008 44276 22060 44285
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 20352 44140 20404 44192
rect 24952 44140 25004 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 6552 43979 6604 43988
rect 6552 43945 6561 43979
rect 6561 43945 6595 43979
rect 6595 43945 6604 43979
rect 6552 43936 6604 43945
rect 7380 43936 7432 43988
rect 8944 43936 8996 43988
rect 17592 43979 17644 43988
rect 17592 43945 17601 43979
rect 17601 43945 17635 43979
rect 17635 43945 17644 43979
rect 17592 43936 17644 43945
rect 19800 43936 19852 43988
rect 9220 43868 9272 43920
rect 16212 43800 16264 43852
rect 18604 43800 18656 43852
rect 20076 43800 20128 43852
rect 10324 43732 10376 43784
rect 10692 43732 10744 43784
rect 11796 43775 11848 43784
rect 11796 43741 11805 43775
rect 11805 43741 11839 43775
rect 11839 43741 11848 43775
rect 11796 43732 11848 43741
rect 8300 43664 8352 43716
rect 10232 43664 10284 43716
rect 10508 43707 10560 43716
rect 10508 43673 10517 43707
rect 10517 43673 10551 43707
rect 10551 43673 10560 43707
rect 10508 43664 10560 43673
rect 12348 43664 12400 43716
rect 9956 43596 10008 43648
rect 13820 43732 13872 43784
rect 15292 43732 15344 43784
rect 15844 43775 15896 43784
rect 15844 43741 15853 43775
rect 15853 43741 15887 43775
rect 15887 43741 15896 43775
rect 15844 43732 15896 43741
rect 18788 43732 18840 43784
rect 16580 43664 16632 43716
rect 20996 43664 21048 43716
rect 13544 43639 13596 43648
rect 13544 43605 13553 43639
rect 13553 43605 13587 43639
rect 13587 43605 13596 43639
rect 13544 43596 13596 43605
rect 17500 43596 17552 43648
rect 25136 43800 25188 43852
rect 22008 43732 22060 43784
rect 24768 43732 24820 43784
rect 23848 43664 23900 43716
rect 22192 43596 22244 43648
rect 22284 43596 22336 43648
rect 25504 43596 25556 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 5540 43435 5592 43444
rect 5540 43401 5549 43435
rect 5549 43401 5583 43435
rect 5583 43401 5592 43435
rect 5540 43392 5592 43401
rect 5172 43256 5224 43308
rect 10692 43392 10744 43444
rect 12164 43392 12216 43444
rect 17224 43392 17276 43444
rect 22192 43392 22244 43444
rect 9496 43324 9548 43376
rect 23848 43324 23900 43376
rect 15200 43256 15252 43308
rect 17500 43256 17552 43308
rect 17684 43256 17736 43308
rect 24860 43256 24912 43308
rect 10048 43188 10100 43240
rect 9496 43052 9548 43104
rect 9956 43052 10008 43104
rect 10416 43052 10468 43104
rect 12348 43120 12400 43172
rect 17408 43231 17460 43240
rect 17408 43197 17417 43231
rect 17417 43197 17451 43231
rect 17451 43197 17460 43231
rect 17408 43188 17460 43197
rect 22008 43231 22060 43240
rect 22008 43197 22017 43231
rect 22017 43197 22051 43231
rect 22051 43197 22060 43231
rect 22008 43188 22060 43197
rect 22652 43188 22704 43240
rect 23756 43188 23808 43240
rect 15384 43052 15436 43104
rect 16672 43052 16724 43104
rect 22100 43052 22152 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 13820 42848 13872 42900
rect 15108 42848 15160 42900
rect 20352 42848 20404 42900
rect 20996 42848 21048 42900
rect 23848 42848 23900 42900
rect 3700 42712 3752 42764
rect 6460 42712 6512 42764
rect 10232 42780 10284 42832
rect 5356 42644 5408 42696
rect 12624 42755 12676 42764
rect 12624 42721 12633 42755
rect 12633 42721 12667 42755
rect 12667 42721 12676 42755
rect 12624 42712 12676 42721
rect 14280 42755 14332 42764
rect 14280 42721 14289 42755
rect 14289 42721 14323 42755
rect 14323 42721 14332 42755
rect 14280 42712 14332 42721
rect 17868 42712 17920 42764
rect 18604 42780 18656 42832
rect 19432 42755 19484 42764
rect 19432 42721 19441 42755
rect 19441 42721 19475 42755
rect 19475 42721 19484 42755
rect 19432 42712 19484 42721
rect 21272 42712 21324 42764
rect 22008 42712 22060 42764
rect 7104 42644 7156 42696
rect 4160 42576 4212 42628
rect 6460 42576 6512 42628
rect 6920 42576 6972 42628
rect 9864 42644 9916 42696
rect 11796 42644 11848 42696
rect 25320 42687 25372 42696
rect 25320 42653 25329 42687
rect 25329 42653 25363 42687
rect 25363 42653 25372 42687
rect 25320 42644 25372 42653
rect 8576 42576 8628 42628
rect 7012 42551 7064 42560
rect 7012 42517 7021 42551
rect 7021 42517 7055 42551
rect 7055 42517 7064 42551
rect 7012 42508 7064 42517
rect 9312 42508 9364 42560
rect 10048 42576 10100 42628
rect 11520 42576 11572 42628
rect 14280 42576 14332 42628
rect 9956 42508 10008 42560
rect 10140 42508 10192 42560
rect 10600 42508 10652 42560
rect 16764 42576 16816 42628
rect 20996 42576 21048 42628
rect 22560 42619 22612 42628
rect 22560 42585 22569 42619
rect 22569 42585 22603 42619
rect 22603 42585 22612 42619
rect 22560 42576 22612 42585
rect 23848 42576 23900 42628
rect 24584 42576 24636 42628
rect 16028 42551 16080 42560
rect 16028 42517 16037 42551
rect 16037 42517 16071 42551
rect 16071 42517 16080 42551
rect 16028 42508 16080 42517
rect 17500 42551 17552 42560
rect 17500 42517 17509 42551
rect 17509 42517 17543 42551
rect 17543 42517 17552 42551
rect 17500 42508 17552 42517
rect 17776 42508 17828 42560
rect 21180 42551 21232 42560
rect 21180 42517 21189 42551
rect 21189 42517 21223 42551
rect 21223 42517 21232 42551
rect 21180 42508 21232 42517
rect 23572 42508 23624 42560
rect 25228 42508 25280 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 1768 42304 1820 42356
rect 8392 42236 8444 42288
rect 9496 42304 9548 42356
rect 11612 42304 11664 42356
rect 19524 42304 19576 42356
rect 20444 42304 20496 42356
rect 22468 42347 22520 42356
rect 22468 42313 22477 42347
rect 22477 42313 22511 42347
rect 22511 42313 22520 42347
rect 22468 42304 22520 42313
rect 12256 42236 12308 42288
rect 14372 42236 14424 42288
rect 18604 42236 18656 42288
rect 21272 42279 21324 42288
rect 21272 42245 21281 42279
rect 21281 42245 21315 42279
rect 21315 42245 21324 42279
rect 21272 42236 21324 42245
rect 22008 42236 22060 42288
rect 3792 42211 3844 42220
rect 3792 42177 3801 42211
rect 3801 42177 3835 42211
rect 3835 42177 3844 42211
rect 3792 42168 3844 42177
rect 11888 42168 11940 42220
rect 15292 42168 15344 42220
rect 17868 42211 17920 42220
rect 17868 42177 17877 42211
rect 17877 42177 17911 42211
rect 17911 42177 17920 42211
rect 17868 42168 17920 42177
rect 19432 42168 19484 42220
rect 20720 42168 20772 42220
rect 23572 42279 23624 42288
rect 23572 42245 23581 42279
rect 23581 42245 23615 42279
rect 23615 42245 23624 42279
rect 23572 42236 23624 42245
rect 24584 42236 24636 42288
rect 8484 42100 8536 42152
rect 11152 42032 11204 42084
rect 13360 42100 13412 42152
rect 16028 42100 16080 42152
rect 18604 42100 18656 42152
rect 19340 42100 19392 42152
rect 21272 42100 21324 42152
rect 21916 42100 21968 42152
rect 22192 42100 22244 42152
rect 9404 41964 9456 42016
rect 11428 41964 11480 42016
rect 13912 41964 13964 42016
rect 14924 41964 14976 42016
rect 21916 41964 21968 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 3424 41760 3476 41812
rect 7840 41803 7892 41812
rect 7840 41769 7849 41803
rect 7849 41769 7883 41803
rect 7883 41769 7892 41803
rect 7840 41760 7892 41769
rect 17224 41760 17276 41812
rect 5632 41692 5684 41744
rect 19064 41692 19116 41744
rect 8484 41667 8536 41676
rect 8484 41633 8493 41667
rect 8493 41633 8527 41667
rect 8527 41633 8536 41667
rect 8484 41624 8536 41633
rect 11704 41624 11756 41676
rect 13360 41624 13412 41676
rect 15292 41667 15344 41676
rect 15292 41633 15301 41667
rect 15301 41633 15335 41667
rect 15335 41633 15344 41667
rect 15292 41624 15344 41633
rect 17868 41624 17920 41676
rect 18788 41624 18840 41676
rect 19708 41624 19760 41676
rect 20260 41692 20312 41744
rect 24952 41692 25004 41744
rect 21180 41624 21232 41676
rect 21732 41624 21784 41676
rect 6276 41556 6328 41608
rect 8300 41556 8352 41608
rect 10600 41556 10652 41608
rect 19432 41556 19484 41608
rect 21088 41556 21140 41608
rect 21824 41556 21876 41608
rect 22744 41556 22796 41608
rect 23204 41599 23256 41608
rect 23204 41565 23213 41599
rect 23213 41565 23247 41599
rect 23247 41565 23256 41599
rect 23204 41556 23256 41565
rect 23940 41556 23992 41608
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 3976 41488 4028 41540
rect 5356 41531 5408 41540
rect 5356 41497 5365 41531
rect 5365 41497 5399 41531
rect 5399 41497 5408 41531
rect 5356 41488 5408 41497
rect 12072 41488 12124 41540
rect 7840 41420 7892 41472
rect 9588 41420 9640 41472
rect 11428 41420 11480 41472
rect 12624 41420 12676 41472
rect 14372 41420 14424 41472
rect 16580 41420 16632 41472
rect 18512 41488 18564 41540
rect 18328 41420 18380 41472
rect 19340 41420 19392 41472
rect 19524 41420 19576 41472
rect 21548 41463 21600 41472
rect 21548 41429 21557 41463
rect 21557 41429 21591 41463
rect 21591 41429 21600 41463
rect 21548 41420 21600 41429
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 3516 41216 3568 41268
rect 7012 41216 7064 41268
rect 7564 41216 7616 41268
rect 8484 41216 8536 41268
rect 11980 41216 12032 41268
rect 12072 41216 12124 41268
rect 15108 41216 15160 41268
rect 17316 41259 17368 41268
rect 17316 41225 17325 41259
rect 17325 41225 17359 41259
rect 17359 41225 17368 41259
rect 17316 41216 17368 41225
rect 13912 41148 13964 41200
rect 14280 41148 14332 41200
rect 20812 41216 20864 41268
rect 21456 41216 21508 41268
rect 22836 41216 22888 41268
rect 4068 41080 4120 41132
rect 8300 41080 8352 41132
rect 12072 41123 12124 41132
rect 12072 41089 12081 41123
rect 12081 41089 12115 41123
rect 12115 41089 12124 41123
rect 12072 41080 12124 41089
rect 13360 41123 13412 41132
rect 13360 41089 13369 41123
rect 13369 41089 13403 41123
rect 13403 41089 13412 41123
rect 13360 41080 13412 41089
rect 18788 41148 18840 41200
rect 19248 41148 19300 41200
rect 21088 41148 21140 41200
rect 22008 41148 22060 41200
rect 22100 41080 22152 41132
rect 23480 41191 23532 41200
rect 23480 41157 23489 41191
rect 23489 41157 23523 41191
rect 23523 41157 23532 41191
rect 23480 41148 23532 41157
rect 24492 41148 24544 41200
rect 6276 41012 6328 41064
rect 7564 41012 7616 41064
rect 9404 41055 9456 41064
rect 9404 41021 9413 41055
rect 9413 41021 9447 41055
rect 9447 41021 9456 41055
rect 9404 41012 9456 41021
rect 11612 41012 11664 41064
rect 12348 41055 12400 41064
rect 12348 41021 12357 41055
rect 12357 41021 12391 41055
rect 12391 41021 12400 41055
rect 12348 41012 12400 41021
rect 14004 41012 14056 41064
rect 18696 41055 18748 41064
rect 18696 41021 18705 41055
rect 18705 41021 18739 41055
rect 18739 41021 18748 41055
rect 18696 41012 18748 41021
rect 19064 41012 19116 41064
rect 22560 41012 22612 41064
rect 11152 40919 11204 40928
rect 11152 40885 11161 40919
rect 11161 40885 11195 40919
rect 11195 40885 11204 40919
rect 11152 40876 11204 40885
rect 14924 40876 14976 40928
rect 16856 40919 16908 40928
rect 16856 40885 16865 40919
rect 16865 40885 16899 40919
rect 16899 40885 16908 40919
rect 16856 40876 16908 40885
rect 18512 40876 18564 40928
rect 18788 40876 18840 40928
rect 19248 40876 19300 40928
rect 20076 40876 20128 40928
rect 21456 40919 21508 40928
rect 21456 40885 21465 40919
rect 21465 40885 21499 40919
rect 21499 40885 21508 40919
rect 21456 40876 21508 40885
rect 23664 40876 23716 40928
rect 25044 40876 25096 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 1584 40672 1636 40724
rect 15200 40672 15252 40724
rect 17684 40672 17736 40724
rect 17868 40672 17920 40724
rect 13820 40604 13872 40656
rect 19064 40604 19116 40656
rect 12164 40536 12216 40588
rect 6276 40511 6328 40520
rect 6276 40477 6285 40511
rect 6285 40477 6319 40511
rect 6319 40477 6328 40511
rect 6276 40468 6328 40477
rect 12624 40536 12676 40588
rect 16396 40579 16448 40588
rect 16396 40545 16405 40579
rect 16405 40545 16439 40579
rect 16439 40545 16448 40579
rect 16396 40536 16448 40545
rect 16488 40536 16540 40588
rect 18604 40536 18656 40588
rect 19616 40536 19668 40588
rect 13452 40468 13504 40520
rect 16672 40468 16724 40520
rect 18328 40468 18380 40520
rect 18512 40468 18564 40520
rect 5080 40400 5132 40452
rect 6552 40443 6604 40452
rect 6552 40409 6561 40443
rect 6561 40409 6595 40443
rect 6595 40409 6604 40443
rect 6552 40400 6604 40409
rect 8300 40400 8352 40452
rect 11428 40443 11480 40452
rect 11428 40409 11437 40443
rect 11437 40409 11471 40443
rect 11471 40409 11480 40443
rect 11428 40400 11480 40409
rect 11796 40400 11848 40452
rect 12164 40443 12216 40452
rect 12164 40409 12173 40443
rect 12173 40409 12207 40443
rect 12207 40409 12216 40443
rect 12164 40400 12216 40409
rect 12348 40400 12400 40452
rect 14280 40400 14332 40452
rect 18604 40400 18656 40452
rect 21364 40672 21416 40724
rect 21088 40579 21140 40588
rect 21088 40545 21097 40579
rect 21097 40545 21131 40579
rect 21131 40545 21140 40579
rect 21088 40536 21140 40545
rect 23572 40536 23624 40588
rect 23664 40468 23716 40520
rect 24952 40468 25004 40520
rect 21272 40400 21324 40452
rect 24400 40400 24452 40452
rect 7564 40332 7616 40384
rect 15752 40332 15804 40384
rect 16212 40375 16264 40384
rect 16212 40341 16221 40375
rect 16221 40341 16255 40375
rect 16255 40341 16264 40375
rect 16212 40332 16264 40341
rect 17684 40375 17736 40384
rect 17684 40341 17693 40375
rect 17693 40341 17727 40375
rect 17727 40341 17736 40375
rect 17684 40332 17736 40341
rect 18328 40332 18380 40384
rect 19708 40332 19760 40384
rect 22836 40375 22888 40384
rect 22836 40341 22845 40375
rect 22845 40341 22879 40375
rect 22879 40341 22888 40375
rect 22836 40332 22888 40341
rect 23572 40332 23624 40384
rect 23664 40375 23716 40384
rect 23664 40341 23673 40375
rect 23673 40341 23707 40375
rect 23707 40341 23716 40375
rect 23664 40332 23716 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 8760 40128 8812 40180
rect 6092 40060 6144 40112
rect 11428 40128 11480 40180
rect 3884 39992 3936 40044
rect 9404 40060 9456 40112
rect 9864 39992 9916 40044
rect 12532 40128 12584 40180
rect 12440 40060 12492 40112
rect 13912 40060 13964 40112
rect 14280 40060 14332 40112
rect 20260 40060 20312 40112
rect 21456 40128 21508 40180
rect 23848 40128 23900 40180
rect 21916 39992 21968 40044
rect 24860 39992 24912 40044
rect 7288 39856 7340 39908
rect 12164 39967 12216 39976
rect 12164 39933 12173 39967
rect 12173 39933 12207 39967
rect 12207 39933 12216 39967
rect 12164 39924 12216 39933
rect 12440 39967 12492 39976
rect 12440 39933 12449 39967
rect 12449 39933 12483 39967
rect 12483 39933 12492 39967
rect 12440 39924 12492 39933
rect 12532 39924 12584 39976
rect 15016 39924 15068 39976
rect 9864 39856 9916 39908
rect 11704 39856 11756 39908
rect 13544 39856 13596 39908
rect 17868 39924 17920 39976
rect 19616 39924 19668 39976
rect 21180 39967 21232 39976
rect 21180 39933 21189 39967
rect 21189 39933 21223 39967
rect 21223 39933 21232 39967
rect 21180 39924 21232 39933
rect 22192 39924 22244 39976
rect 22284 39924 22336 39976
rect 16580 39856 16632 39908
rect 6552 39788 6604 39840
rect 11244 39788 11296 39840
rect 11612 39788 11664 39840
rect 13912 39831 13964 39840
rect 13912 39797 13921 39831
rect 13921 39797 13955 39831
rect 13955 39797 13964 39831
rect 13912 39788 13964 39797
rect 14004 39788 14056 39840
rect 15200 39831 15252 39840
rect 15200 39797 15209 39831
rect 15209 39797 15243 39831
rect 15243 39797 15252 39831
rect 15200 39788 15252 39797
rect 17500 39788 17552 39840
rect 18052 39788 18104 39840
rect 18420 39788 18472 39840
rect 18788 39788 18840 39840
rect 20536 39856 20588 39908
rect 25136 39856 25188 39908
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 6920 39584 6972 39636
rect 7196 39584 7248 39636
rect 7656 39627 7708 39636
rect 7656 39593 7665 39627
rect 7665 39593 7699 39627
rect 7699 39593 7708 39627
rect 7656 39584 7708 39593
rect 11152 39584 11204 39636
rect 11244 39584 11296 39636
rect 9864 39516 9916 39568
rect 11704 39516 11756 39568
rect 6920 39448 6972 39500
rect 9036 39448 9088 39500
rect 12164 39448 12216 39500
rect 12440 39448 12492 39500
rect 13636 39584 13688 39636
rect 16396 39584 16448 39636
rect 18788 39584 18840 39636
rect 19524 39627 19576 39636
rect 19524 39593 19533 39627
rect 19533 39593 19567 39627
rect 19567 39593 19576 39627
rect 19524 39584 19576 39593
rect 20720 39627 20772 39636
rect 20720 39593 20729 39627
rect 20729 39593 20763 39627
rect 20763 39593 20772 39627
rect 20720 39584 20772 39593
rect 23664 39584 23716 39636
rect 7472 39380 7524 39432
rect 9496 39423 9548 39432
rect 9496 39389 9505 39423
rect 9505 39389 9539 39423
rect 9539 39389 9548 39423
rect 9496 39380 9548 39389
rect 12348 39380 12400 39432
rect 12532 39380 12584 39432
rect 12716 39380 12768 39432
rect 13912 39448 13964 39500
rect 16396 39491 16448 39500
rect 16396 39457 16405 39491
rect 16405 39457 16439 39491
rect 16439 39457 16448 39491
rect 16396 39448 16448 39457
rect 13544 39380 13596 39432
rect 15200 39380 15252 39432
rect 19248 39516 19300 39568
rect 21824 39516 21876 39568
rect 25780 39516 25832 39568
rect 9680 39312 9732 39364
rect 12256 39312 12308 39364
rect 7656 39244 7708 39296
rect 9404 39244 9456 39296
rect 12164 39244 12216 39296
rect 12348 39244 12400 39296
rect 12992 39287 13044 39296
rect 12992 39253 13001 39287
rect 13001 39253 13035 39287
rect 13035 39253 13044 39287
rect 12992 39244 13044 39253
rect 17408 39380 17460 39432
rect 15568 39244 15620 39296
rect 17592 39448 17644 39500
rect 18052 39448 18104 39500
rect 20352 39448 20404 39500
rect 21088 39448 21140 39500
rect 21640 39448 21692 39500
rect 17592 39312 17644 39364
rect 17960 39312 18012 39364
rect 19616 39312 19668 39364
rect 18972 39244 19024 39296
rect 19892 39287 19944 39296
rect 19892 39253 19901 39287
rect 19901 39253 19935 39287
rect 19935 39253 19944 39287
rect 19892 39244 19944 39253
rect 21824 39312 21876 39364
rect 22192 39380 22244 39432
rect 22836 39448 22888 39500
rect 25044 39448 25096 39500
rect 24032 39423 24084 39432
rect 24032 39389 24041 39423
rect 24041 39389 24075 39423
rect 24075 39389 24084 39423
rect 24032 39380 24084 39389
rect 24952 39423 25004 39432
rect 24952 39389 24961 39423
rect 24961 39389 24995 39423
rect 24995 39389 25004 39423
rect 24952 39380 25004 39389
rect 22468 39312 22520 39364
rect 25412 39312 25464 39364
rect 20628 39244 20680 39296
rect 21916 39287 21968 39296
rect 21916 39253 21925 39287
rect 21925 39253 21959 39287
rect 21959 39253 21968 39287
rect 21916 39244 21968 39253
rect 22284 39287 22336 39296
rect 22284 39253 22293 39287
rect 22293 39253 22327 39287
rect 22327 39253 22336 39287
rect 22284 39244 22336 39253
rect 24308 39244 24360 39296
rect 25044 39287 25096 39296
rect 25044 39253 25053 39287
rect 25053 39253 25087 39287
rect 25087 39253 25096 39287
rect 25044 39244 25096 39253
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 9772 39040 9824 39092
rect 11888 39040 11940 39092
rect 14004 39083 14056 39092
rect 14004 39049 14013 39083
rect 14013 39049 14047 39083
rect 14047 39049 14056 39083
rect 14004 39040 14056 39049
rect 16856 39040 16908 39092
rect 12716 38972 12768 39024
rect 12992 38972 13044 39024
rect 16580 38972 16632 39024
rect 17316 38972 17368 39024
rect 18604 39040 18656 39092
rect 18420 38972 18472 39024
rect 19708 39040 19760 39092
rect 22376 39040 22428 39092
rect 940 38904 992 38956
rect 10048 38947 10100 38956
rect 10048 38913 10057 38947
rect 10057 38913 10091 38947
rect 10091 38913 10100 38947
rect 10048 38904 10100 38913
rect 15844 38947 15896 38956
rect 15844 38913 15853 38947
rect 15853 38913 15887 38947
rect 15887 38913 15896 38947
rect 15844 38904 15896 38913
rect 21088 38972 21140 39024
rect 22744 38972 22796 39024
rect 24400 38972 24452 39024
rect 9312 38836 9364 38888
rect 12256 38879 12308 38888
rect 12256 38845 12265 38879
rect 12265 38845 12299 38879
rect 12299 38845 12308 38879
rect 12256 38836 12308 38845
rect 9496 38768 9548 38820
rect 1860 38700 1912 38752
rect 8668 38743 8720 38752
rect 8668 38709 8677 38743
rect 8677 38709 8711 38743
rect 8711 38709 8720 38743
rect 8668 38700 8720 38709
rect 11152 38700 11204 38752
rect 11612 38768 11664 38820
rect 13820 38836 13872 38888
rect 14556 38836 14608 38888
rect 16028 38879 16080 38888
rect 16028 38845 16037 38879
rect 16037 38845 16071 38879
rect 16071 38845 16080 38879
rect 16028 38836 16080 38845
rect 17040 38836 17092 38888
rect 16212 38768 16264 38820
rect 13360 38700 13412 38752
rect 16488 38700 16540 38752
rect 16672 38700 16724 38752
rect 20444 38879 20496 38888
rect 20444 38845 20453 38879
rect 20453 38845 20487 38879
rect 20487 38845 20496 38879
rect 20444 38836 20496 38845
rect 19616 38768 19668 38820
rect 22836 38904 22888 38956
rect 23388 38879 23440 38888
rect 23388 38845 23397 38879
rect 23397 38845 23431 38879
rect 23431 38845 23440 38879
rect 23388 38836 23440 38845
rect 24216 38836 24268 38888
rect 19524 38700 19576 38752
rect 22008 38743 22060 38752
rect 22008 38709 22017 38743
rect 22017 38709 22051 38743
rect 22051 38709 22060 38743
rect 22008 38700 22060 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 6920 38496 6972 38548
rect 7564 38496 7616 38548
rect 7840 38539 7892 38548
rect 7840 38505 7849 38539
rect 7849 38505 7883 38539
rect 7883 38505 7892 38539
rect 7840 38496 7892 38505
rect 9404 38496 9456 38548
rect 11520 38496 11572 38548
rect 6276 38360 6328 38412
rect 7564 38360 7616 38412
rect 11244 38428 11296 38480
rect 7380 38292 7432 38344
rect 8024 38292 8076 38344
rect 8668 38292 8720 38344
rect 5540 38224 5592 38276
rect 10324 38360 10376 38412
rect 11336 38403 11388 38412
rect 11336 38369 11345 38403
rect 11345 38369 11379 38403
rect 11379 38369 11388 38403
rect 11336 38360 11388 38369
rect 9588 38292 9640 38344
rect 12164 38428 12216 38480
rect 16764 38539 16816 38548
rect 16764 38505 16773 38539
rect 16773 38505 16807 38539
rect 16807 38505 16816 38539
rect 16764 38496 16816 38505
rect 22284 38496 22336 38548
rect 22560 38496 22612 38548
rect 23480 38496 23532 38548
rect 12348 38360 12400 38412
rect 13360 38360 13412 38412
rect 9772 38224 9824 38276
rect 7840 38156 7892 38208
rect 8024 38156 8076 38208
rect 8392 38156 8444 38208
rect 11336 38224 11388 38276
rect 14556 38292 14608 38344
rect 16304 38403 16356 38412
rect 16304 38369 16313 38403
rect 16313 38369 16347 38403
rect 16347 38369 16356 38403
rect 16304 38360 16356 38369
rect 17224 38403 17276 38412
rect 17224 38369 17233 38403
rect 17233 38369 17267 38403
rect 17267 38369 17276 38403
rect 17224 38360 17276 38369
rect 22100 38428 22152 38480
rect 19340 38360 19392 38412
rect 20076 38403 20128 38412
rect 20076 38369 20085 38403
rect 20085 38369 20119 38403
rect 20119 38369 20128 38403
rect 20076 38360 20128 38369
rect 21272 38403 21324 38412
rect 21272 38369 21281 38403
rect 21281 38369 21315 38403
rect 21315 38369 21324 38403
rect 21272 38360 21324 38369
rect 25688 38428 25740 38480
rect 22560 38360 22612 38412
rect 23296 38360 23348 38412
rect 11060 38199 11112 38208
rect 11060 38165 11069 38199
rect 11069 38165 11103 38199
rect 11103 38165 11112 38199
rect 11060 38156 11112 38165
rect 11244 38156 11296 38208
rect 12348 38199 12400 38208
rect 12348 38165 12357 38199
rect 12357 38165 12391 38199
rect 12391 38165 12400 38199
rect 12348 38156 12400 38165
rect 14372 38199 14424 38208
rect 14372 38165 14381 38199
rect 14381 38165 14415 38199
rect 14415 38165 14424 38199
rect 14372 38156 14424 38165
rect 15660 38199 15712 38208
rect 15660 38165 15669 38199
rect 15669 38165 15703 38199
rect 15703 38165 15712 38199
rect 15660 38156 15712 38165
rect 17592 38224 17644 38276
rect 18604 38224 18656 38276
rect 19984 38224 20036 38276
rect 21548 38292 21600 38344
rect 25412 38292 25464 38344
rect 21456 38224 21508 38276
rect 16120 38199 16172 38208
rect 16120 38165 16129 38199
rect 16129 38165 16163 38199
rect 16163 38165 16172 38199
rect 16120 38156 16172 38165
rect 16212 38199 16264 38208
rect 16212 38165 16221 38199
rect 16221 38165 16255 38199
rect 16255 38165 16264 38199
rect 16212 38156 16264 38165
rect 17132 38199 17184 38208
rect 17132 38165 17141 38199
rect 17141 38165 17175 38199
rect 17175 38165 17184 38199
rect 17132 38156 17184 38165
rect 20260 38156 20312 38208
rect 20720 38156 20772 38208
rect 21824 38156 21876 38208
rect 22468 38156 22520 38208
rect 23664 38156 23716 38208
rect 25136 38199 25188 38208
rect 25136 38165 25145 38199
rect 25145 38165 25179 38199
rect 25179 38165 25188 38199
rect 25136 38156 25188 38165
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 6552 37952 6604 38004
rect 7012 37952 7064 38004
rect 10324 37952 10376 38004
rect 11152 37952 11204 38004
rect 11336 37952 11388 38004
rect 12808 37952 12860 38004
rect 15844 37952 15896 38004
rect 5540 37884 5592 37936
rect 8300 37884 8352 37936
rect 14188 37884 14240 37936
rect 16580 37884 16632 37936
rect 18788 37995 18840 38004
rect 18788 37961 18797 37995
rect 18797 37961 18831 37995
rect 18831 37961 18840 37995
rect 18788 37952 18840 37961
rect 19616 37952 19668 38004
rect 22376 37952 22428 38004
rect 22744 37952 22796 38004
rect 23756 37952 23808 38004
rect 24216 37952 24268 38004
rect 19432 37884 19484 37936
rect 23296 37884 23348 37936
rect 24492 37884 24544 37936
rect 7564 37859 7616 37868
rect 7564 37825 7573 37859
rect 7573 37825 7607 37859
rect 7607 37825 7616 37859
rect 7564 37816 7616 37825
rect 10232 37816 10284 37868
rect 11060 37816 11112 37868
rect 15292 37859 15344 37868
rect 15292 37825 15301 37859
rect 15301 37825 15335 37859
rect 15335 37825 15344 37859
rect 15292 37816 15344 37825
rect 16120 37816 16172 37868
rect 18420 37816 18472 37868
rect 19064 37816 19116 37868
rect 4528 37791 4580 37800
rect 4528 37757 4537 37791
rect 4537 37757 4571 37791
rect 4571 37757 4580 37791
rect 4528 37748 4580 37757
rect 9312 37748 9364 37800
rect 9036 37680 9088 37732
rect 10600 37791 10652 37800
rect 10600 37757 10609 37791
rect 10609 37757 10643 37791
rect 10643 37757 10652 37791
rect 10600 37748 10652 37757
rect 10692 37791 10744 37800
rect 10692 37757 10701 37791
rect 10701 37757 10735 37791
rect 10735 37757 10744 37791
rect 10692 37748 10744 37757
rect 11520 37748 11572 37800
rect 12072 37680 12124 37732
rect 14188 37748 14240 37800
rect 14924 37748 14976 37800
rect 17040 37791 17092 37800
rect 17040 37757 17049 37791
rect 17049 37757 17083 37791
rect 17083 37757 17092 37791
rect 17040 37748 17092 37757
rect 17868 37748 17920 37800
rect 13820 37680 13872 37732
rect 4988 37612 5040 37664
rect 11060 37612 11112 37664
rect 12164 37612 12216 37664
rect 12808 37612 12860 37664
rect 16764 37680 16816 37732
rect 20536 37680 20588 37732
rect 22652 37748 22704 37800
rect 23388 37748 23440 37800
rect 14924 37655 14976 37664
rect 14924 37621 14933 37655
rect 14933 37621 14967 37655
rect 14967 37621 14976 37655
rect 14924 37612 14976 37621
rect 18052 37612 18104 37664
rect 18512 37612 18564 37664
rect 19616 37655 19668 37664
rect 19616 37621 19625 37655
rect 19625 37621 19659 37655
rect 19659 37621 19668 37655
rect 19616 37612 19668 37621
rect 20996 37612 21048 37664
rect 21548 37612 21600 37664
rect 25228 37612 25280 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 6184 37408 6236 37460
rect 7012 37408 7064 37460
rect 10692 37408 10744 37460
rect 8392 37340 8444 37392
rect 11520 37340 11572 37392
rect 15384 37340 15436 37392
rect 15660 37408 15712 37460
rect 22376 37408 22428 37460
rect 22744 37408 22796 37460
rect 16396 37340 16448 37392
rect 6920 37272 6972 37324
rect 7012 37272 7064 37324
rect 10324 37315 10376 37324
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 10416 37272 10468 37324
rect 16212 37272 16264 37324
rect 4988 37204 5040 37256
rect 7288 37247 7340 37256
rect 7288 37213 7297 37247
rect 7297 37213 7331 37247
rect 7331 37213 7340 37247
rect 7288 37204 7340 37213
rect 8760 37204 8812 37256
rect 5540 37136 5592 37188
rect 9864 37136 9916 37188
rect 7748 37111 7800 37120
rect 7748 37077 7757 37111
rect 7757 37077 7791 37111
rect 7791 37077 7800 37111
rect 7748 37068 7800 37077
rect 10140 37111 10192 37120
rect 10140 37077 10149 37111
rect 10149 37077 10183 37111
rect 10183 37077 10192 37111
rect 10140 37068 10192 37077
rect 10232 37068 10284 37120
rect 13636 37204 13688 37256
rect 17224 37340 17276 37392
rect 18052 37272 18104 37324
rect 19340 37340 19392 37392
rect 21088 37272 21140 37324
rect 21640 37315 21692 37324
rect 21640 37281 21649 37315
rect 21649 37281 21683 37315
rect 21683 37281 21692 37315
rect 21640 37272 21692 37281
rect 22192 37272 22244 37324
rect 19616 37204 19668 37256
rect 15292 37136 15344 37188
rect 19432 37179 19484 37188
rect 19432 37145 19441 37179
rect 19441 37145 19475 37179
rect 19475 37145 19484 37179
rect 19432 37136 19484 37145
rect 20168 37179 20220 37188
rect 20168 37145 20177 37179
rect 20177 37145 20211 37179
rect 20211 37145 20220 37179
rect 20168 37136 20220 37145
rect 11336 37111 11388 37120
rect 11336 37077 11345 37111
rect 11345 37077 11379 37111
rect 11379 37077 11388 37111
rect 11336 37068 11388 37077
rect 15476 37111 15528 37120
rect 15476 37077 15485 37111
rect 15485 37077 15519 37111
rect 15519 37077 15528 37111
rect 15476 37068 15528 37077
rect 16672 37068 16724 37120
rect 16948 37068 17000 37120
rect 17592 37111 17644 37120
rect 17592 37077 17601 37111
rect 17601 37077 17635 37111
rect 17635 37077 17644 37111
rect 17592 37068 17644 37077
rect 21180 37068 21232 37120
rect 22928 37136 22980 37188
rect 23756 37247 23808 37256
rect 23756 37213 23765 37247
rect 23765 37213 23799 37247
rect 23799 37213 23808 37247
rect 23756 37204 23808 37213
rect 24860 37204 24912 37256
rect 24492 37136 24544 37188
rect 22652 37068 22704 37120
rect 23112 37111 23164 37120
rect 23112 37077 23121 37111
rect 23121 37077 23155 37111
rect 23155 37077 23164 37111
rect 23112 37068 23164 37077
rect 23388 37068 23440 37120
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 5172 36907 5224 36916
rect 5172 36873 5181 36907
rect 5181 36873 5215 36907
rect 5215 36873 5224 36907
rect 5172 36864 5224 36873
rect 9128 36864 9180 36916
rect 9312 36907 9364 36916
rect 9312 36873 9321 36907
rect 9321 36873 9355 36907
rect 9355 36873 9364 36907
rect 9312 36864 9364 36873
rect 10140 36864 10192 36916
rect 6828 36796 6880 36848
rect 8300 36796 8352 36848
rect 12716 36864 12768 36916
rect 14372 36864 14424 36916
rect 15292 36907 15344 36916
rect 15292 36873 15301 36907
rect 15301 36873 15335 36907
rect 15335 36873 15344 36907
rect 15292 36864 15344 36873
rect 16028 36864 16080 36916
rect 16856 36796 16908 36848
rect 940 36728 992 36780
rect 4620 36728 4672 36780
rect 9312 36728 9364 36780
rect 13544 36728 13596 36780
rect 17132 36728 17184 36780
rect 17500 36728 17552 36780
rect 18328 36864 18380 36916
rect 19248 36864 19300 36916
rect 22008 36864 22060 36916
rect 17684 36796 17736 36848
rect 19800 36796 19852 36848
rect 24584 36864 24636 36916
rect 22560 36796 22612 36848
rect 23112 36796 23164 36848
rect 24492 36796 24544 36848
rect 19432 36728 19484 36780
rect 22284 36728 22336 36780
rect 25320 36771 25372 36780
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 4528 36592 4580 36644
rect 5264 36592 5316 36644
rect 6092 36660 6144 36712
rect 7564 36703 7616 36712
rect 7564 36669 7573 36703
rect 7573 36669 7607 36703
rect 7607 36669 7616 36703
rect 7564 36660 7616 36669
rect 9588 36660 9640 36712
rect 10232 36703 10284 36712
rect 10232 36669 10241 36703
rect 10241 36669 10275 36703
rect 10275 36669 10284 36703
rect 10232 36660 10284 36669
rect 9496 36592 9548 36644
rect 13452 36703 13504 36712
rect 13452 36669 13461 36703
rect 13461 36669 13495 36703
rect 13495 36669 13504 36703
rect 13452 36660 13504 36669
rect 16212 36660 16264 36712
rect 18512 36703 18564 36712
rect 18512 36669 18521 36703
rect 18521 36669 18555 36703
rect 18555 36669 18564 36703
rect 18512 36660 18564 36669
rect 16120 36592 16172 36644
rect 18420 36592 18472 36644
rect 19708 36660 19760 36712
rect 22652 36660 22704 36712
rect 20720 36592 20772 36644
rect 21364 36592 21416 36644
rect 25504 36660 25556 36712
rect 3424 36524 3476 36576
rect 7196 36524 7248 36576
rect 9956 36524 10008 36576
rect 16304 36524 16356 36576
rect 20628 36524 20680 36576
rect 22468 36524 22520 36576
rect 22836 36524 22888 36576
rect 23480 36524 23532 36576
rect 24860 36524 24912 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7840 36363 7892 36372
rect 7840 36329 7849 36363
rect 7849 36329 7883 36363
rect 7883 36329 7892 36363
rect 7840 36320 7892 36329
rect 9036 36320 9088 36372
rect 12532 36320 12584 36372
rect 13084 36320 13136 36372
rect 18604 36320 18656 36372
rect 8576 36252 8628 36304
rect 8760 36252 8812 36304
rect 7564 36184 7616 36236
rect 12716 36184 12768 36236
rect 16764 36252 16816 36304
rect 18696 36252 18748 36304
rect 17684 36227 17736 36236
rect 17684 36193 17693 36227
rect 17693 36193 17727 36227
rect 17727 36193 17736 36227
rect 17684 36184 17736 36193
rect 4988 36116 5040 36168
rect 6092 36159 6144 36168
rect 6092 36125 6101 36159
rect 6101 36125 6135 36159
rect 6135 36125 6144 36159
rect 6092 36116 6144 36125
rect 11428 36116 11480 36168
rect 5540 35980 5592 36032
rect 6828 36048 6880 36100
rect 11796 36091 11848 36100
rect 11796 36057 11805 36091
rect 11805 36057 11839 36091
rect 11839 36057 11848 36091
rect 11796 36048 11848 36057
rect 13360 36116 13412 36168
rect 15200 36116 15252 36168
rect 16304 36159 16356 36168
rect 16304 36125 16313 36159
rect 16313 36125 16347 36159
rect 16347 36125 16356 36159
rect 16304 36116 16356 36125
rect 21456 36363 21508 36372
rect 21456 36329 21465 36363
rect 21465 36329 21499 36363
rect 21499 36329 21508 36363
rect 21456 36320 21508 36329
rect 21916 36320 21968 36372
rect 22744 36320 22796 36372
rect 22836 36320 22888 36372
rect 23756 36320 23808 36372
rect 21272 36252 21324 36304
rect 20628 36227 20680 36236
rect 20628 36193 20637 36227
rect 20637 36193 20671 36227
rect 20671 36193 20680 36227
rect 20628 36184 20680 36193
rect 21732 36184 21784 36236
rect 23480 36184 23532 36236
rect 23664 36184 23716 36236
rect 24216 36184 24268 36236
rect 25044 36116 25096 36168
rect 25504 36116 25556 36168
rect 16028 36048 16080 36100
rect 17592 36091 17644 36100
rect 17592 36057 17601 36091
rect 17601 36057 17635 36091
rect 17635 36057 17644 36091
rect 17592 36048 17644 36057
rect 19064 36048 19116 36100
rect 19248 36048 19300 36100
rect 20352 36091 20404 36100
rect 20352 36057 20361 36091
rect 20361 36057 20395 36091
rect 20395 36057 20404 36091
rect 20352 36048 20404 36057
rect 21180 36048 21232 36100
rect 22008 36048 22060 36100
rect 22100 36048 22152 36100
rect 24124 36048 24176 36100
rect 8300 35980 8352 36032
rect 9680 35980 9732 36032
rect 12440 36023 12492 36032
rect 12440 35989 12449 36023
rect 12449 35989 12483 36023
rect 12483 35989 12492 36023
rect 12440 35980 12492 35989
rect 15292 35980 15344 36032
rect 18512 35980 18564 36032
rect 19340 35980 19392 36032
rect 20720 35980 20772 36032
rect 20812 35980 20864 36032
rect 22376 35980 22428 36032
rect 22836 35980 22888 36032
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 7012 35776 7064 35828
rect 9588 35776 9640 35828
rect 5540 35708 5592 35760
rect 9680 35708 9732 35760
rect 10140 35708 10192 35760
rect 4160 35436 4212 35488
rect 6828 35572 6880 35624
rect 9220 35572 9272 35624
rect 10692 35572 10744 35624
rect 11060 35572 11112 35624
rect 4988 35436 5040 35488
rect 12808 35776 12860 35828
rect 13636 35776 13688 35828
rect 15108 35776 15160 35828
rect 16856 35819 16908 35828
rect 16856 35785 16865 35819
rect 16865 35785 16899 35819
rect 16899 35785 16908 35819
rect 16856 35776 16908 35785
rect 18604 35776 18656 35828
rect 17040 35708 17092 35760
rect 20168 35776 20220 35828
rect 13360 35640 13412 35692
rect 11796 35615 11848 35624
rect 11796 35581 11805 35615
rect 11805 35581 11839 35615
rect 11839 35581 11848 35615
rect 11796 35572 11848 35581
rect 14188 35572 14240 35624
rect 13084 35504 13136 35556
rect 16304 35640 16356 35692
rect 18788 35708 18840 35760
rect 19340 35708 19392 35760
rect 23480 35751 23532 35760
rect 23480 35717 23489 35751
rect 23489 35717 23523 35751
rect 23523 35717 23532 35751
rect 23480 35708 23532 35717
rect 24492 35708 24544 35760
rect 15292 35572 15344 35624
rect 16396 35572 16448 35624
rect 17316 35615 17368 35624
rect 17316 35581 17325 35615
rect 17325 35581 17359 35615
rect 17359 35581 17368 35615
rect 17316 35572 17368 35581
rect 17132 35504 17184 35556
rect 13452 35436 13504 35488
rect 14004 35479 14056 35488
rect 14004 35445 14013 35479
rect 14013 35445 14047 35479
rect 14047 35445 14056 35479
rect 14004 35436 14056 35445
rect 14648 35436 14700 35488
rect 19248 35572 19300 35624
rect 22744 35640 22796 35692
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 22652 35572 22704 35624
rect 19340 35436 19392 35488
rect 21088 35436 21140 35488
rect 22744 35436 22796 35488
rect 23296 35436 23348 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 7104 35232 7156 35284
rect 10048 35232 10100 35284
rect 15568 35232 15620 35284
rect 17316 35232 17368 35284
rect 19708 35232 19760 35284
rect 21548 35232 21600 35284
rect 23664 35232 23716 35284
rect 7288 35164 7340 35216
rect 7564 35164 7616 35216
rect 9220 35164 9272 35216
rect 11796 35164 11848 35216
rect 6920 35096 6972 35148
rect 9588 35096 9640 35148
rect 4988 35028 5040 35080
rect 9956 35071 10008 35080
rect 9956 35037 9965 35071
rect 9965 35037 9999 35071
rect 9999 35037 10008 35071
rect 9956 35028 10008 35037
rect 13452 35164 13504 35216
rect 13360 35028 13412 35080
rect 13636 35096 13688 35148
rect 16580 35096 16632 35148
rect 17132 35164 17184 35216
rect 17960 35164 18012 35216
rect 18972 35164 19024 35216
rect 19340 35164 19392 35216
rect 19616 35096 19668 35148
rect 20720 35096 20772 35148
rect 22100 35096 22152 35148
rect 22468 35096 22520 35148
rect 23204 35096 23256 35148
rect 23296 35096 23348 35148
rect 13820 35028 13872 35080
rect 14832 35028 14884 35080
rect 15200 35071 15252 35080
rect 15200 35037 15209 35071
rect 15209 35037 15243 35071
rect 15243 35037 15252 35071
rect 15200 35028 15252 35037
rect 25136 35028 25188 35080
rect 25412 35028 25464 35080
rect 5540 34960 5592 35012
rect 6828 34960 6880 35012
rect 10324 34960 10376 35012
rect 7840 34892 7892 34944
rect 9588 34892 9640 34944
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 10140 34892 10192 34944
rect 18696 34960 18748 35012
rect 14188 34892 14240 34944
rect 18880 34892 18932 34944
rect 20076 34960 20128 35012
rect 20720 34960 20772 35012
rect 23204 34935 23256 34944
rect 23204 34901 23213 34935
rect 23213 34901 23247 34935
rect 23247 34901 23256 34935
rect 23204 34892 23256 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 3332 34688 3384 34740
rect 4160 34688 4212 34740
rect 5264 34731 5316 34740
rect 5264 34697 5273 34731
rect 5273 34697 5307 34731
rect 5307 34697 5316 34731
rect 5264 34688 5316 34697
rect 6552 34688 6604 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 5540 34620 5592 34672
rect 7012 34663 7064 34672
rect 7012 34629 7021 34663
rect 7021 34629 7055 34663
rect 7055 34629 7064 34663
rect 7012 34620 7064 34629
rect 7656 34688 7708 34740
rect 11980 34688 12032 34740
rect 12072 34688 12124 34740
rect 13360 34620 13412 34672
rect 15016 34620 15068 34672
rect 17040 34620 17092 34672
rect 19064 34620 19116 34672
rect 4160 34348 4212 34400
rect 7656 34484 7708 34536
rect 11704 34595 11756 34604
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 21180 34688 21232 34740
rect 23388 34688 23440 34740
rect 25044 34688 25096 34740
rect 20996 34620 21048 34672
rect 22560 34620 22612 34672
rect 24308 34620 24360 34672
rect 8300 34416 8352 34468
rect 12624 34484 12676 34536
rect 13360 34484 13412 34536
rect 17132 34527 17184 34536
rect 17132 34493 17141 34527
rect 17141 34493 17175 34527
rect 17175 34493 17184 34527
rect 17132 34484 17184 34493
rect 18328 34484 18380 34536
rect 14832 34416 14884 34468
rect 19248 34484 19300 34536
rect 7748 34348 7800 34400
rect 8484 34391 8536 34400
rect 8484 34357 8493 34391
rect 8493 34357 8527 34391
rect 8527 34357 8536 34391
rect 8484 34348 8536 34357
rect 14556 34348 14608 34400
rect 15108 34348 15160 34400
rect 23204 34552 23256 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 19524 34527 19576 34536
rect 19524 34493 19533 34527
rect 19533 34493 19567 34527
rect 19567 34493 19576 34527
rect 19524 34484 19576 34493
rect 21640 34416 21692 34468
rect 22468 34416 22520 34468
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 4160 34144 4212 34196
rect 5356 34144 5408 34196
rect 6736 34144 6788 34196
rect 9128 34187 9180 34196
rect 9128 34153 9137 34187
rect 9137 34153 9171 34187
rect 9171 34153 9180 34187
rect 9128 34144 9180 34153
rect 12256 34144 12308 34196
rect 17132 34144 17184 34196
rect 20996 34144 21048 34196
rect 6828 34008 6880 34060
rect 11704 34076 11756 34128
rect 12348 34076 12400 34128
rect 14740 34076 14792 34128
rect 19892 34076 19944 34128
rect 23296 34076 23348 34128
rect 24860 34076 24912 34128
rect 12256 34008 12308 34060
rect 4896 33983 4948 33992
rect 4896 33949 4905 33983
rect 4905 33949 4939 33983
rect 4939 33949 4948 33983
rect 4896 33940 4948 33949
rect 12348 33940 12400 33992
rect 12532 34051 12584 34060
rect 12532 34017 12541 34051
rect 12541 34017 12575 34051
rect 12575 34017 12584 34051
rect 12532 34008 12584 34017
rect 13452 34008 13504 34060
rect 18420 34008 18472 34060
rect 20536 34008 20588 34060
rect 23572 34008 23624 34060
rect 17040 33940 17092 33992
rect 17960 33940 18012 33992
rect 5632 33872 5684 33924
rect 11888 33872 11940 33924
rect 11980 33804 12032 33856
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 13268 33872 13320 33924
rect 18972 33872 19024 33924
rect 20352 33940 20404 33992
rect 23848 33983 23900 33992
rect 23848 33949 23857 33983
rect 23857 33949 23891 33983
rect 23891 33949 23900 33983
rect 23848 33940 23900 33949
rect 12808 33804 12860 33856
rect 14004 33804 14056 33856
rect 16580 33804 16632 33856
rect 19800 33804 19852 33856
rect 20812 33804 20864 33856
rect 21916 33804 21968 33856
rect 24492 33872 24544 33924
rect 22468 33847 22520 33856
rect 22468 33813 22477 33847
rect 22477 33813 22511 33847
rect 22511 33813 22520 33847
rect 22468 33804 22520 33813
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 7012 33600 7064 33652
rect 8576 33532 8628 33584
rect 9496 33643 9548 33652
rect 9496 33609 9505 33643
rect 9505 33609 9539 33643
rect 9539 33609 9548 33643
rect 9496 33600 9548 33609
rect 9864 33600 9916 33652
rect 10232 33600 10284 33652
rect 12808 33600 12860 33652
rect 13912 33643 13964 33652
rect 13912 33609 13921 33643
rect 13921 33609 13955 33643
rect 13955 33609 13964 33643
rect 13912 33600 13964 33609
rect 14924 33600 14976 33652
rect 20720 33600 20772 33652
rect 20812 33600 20864 33652
rect 23848 33600 23900 33652
rect 14004 33532 14056 33584
rect 14740 33532 14792 33584
rect 17132 33532 17184 33584
rect 23296 33532 23348 33584
rect 23756 33532 23808 33584
rect 24492 33532 24544 33584
rect 7748 33439 7800 33448
rect 7748 33405 7757 33439
rect 7757 33405 7791 33439
rect 7791 33405 7800 33439
rect 7748 33396 7800 33405
rect 9404 33396 9456 33448
rect 10416 33439 10468 33448
rect 10416 33405 10425 33439
rect 10425 33405 10459 33439
rect 10459 33405 10468 33439
rect 10416 33396 10468 33405
rect 15016 33507 15068 33516
rect 15016 33473 15025 33507
rect 15025 33473 15059 33507
rect 15059 33473 15068 33507
rect 15016 33464 15068 33473
rect 15108 33464 15160 33516
rect 10324 33328 10376 33380
rect 11060 33328 11112 33380
rect 13360 33328 13412 33380
rect 14188 33396 14240 33448
rect 10508 33260 10560 33312
rect 12624 33260 12676 33312
rect 13268 33260 13320 33312
rect 13452 33303 13504 33312
rect 13452 33269 13461 33303
rect 13461 33269 13495 33303
rect 13495 33269 13504 33303
rect 13452 33260 13504 33269
rect 13544 33260 13596 33312
rect 18972 33464 19024 33516
rect 19984 33439 20036 33448
rect 19984 33405 19993 33439
rect 19993 33405 20027 33439
rect 20027 33405 20036 33439
rect 19984 33396 20036 33405
rect 21732 33464 21784 33516
rect 20352 33396 20404 33448
rect 22652 33396 22704 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 20168 33328 20220 33380
rect 15108 33260 15160 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 9312 33056 9364 33108
rect 9588 33056 9640 33108
rect 15016 33056 15068 33108
rect 20444 33056 20496 33108
rect 20996 33056 21048 33108
rect 21824 33056 21876 33108
rect 23020 33056 23072 33108
rect 23388 33056 23440 33108
rect 6828 32988 6880 33040
rect 12716 32988 12768 33040
rect 15844 32988 15896 33040
rect 4896 32920 4948 32972
rect 7748 32920 7800 32972
rect 9404 32920 9456 32972
rect 8392 32852 8444 32904
rect 13820 32920 13872 32972
rect 16120 32963 16172 32972
rect 16120 32929 16129 32963
rect 16129 32929 16163 32963
rect 16163 32929 16172 32963
rect 16120 32920 16172 32929
rect 16304 32963 16356 32972
rect 16304 32929 16313 32963
rect 16313 32929 16347 32963
rect 16347 32929 16356 32963
rect 16304 32920 16356 32929
rect 16856 32963 16908 32972
rect 16856 32929 16865 32963
rect 16865 32929 16899 32963
rect 16899 32929 16908 32963
rect 16856 32920 16908 32929
rect 18972 32988 19024 33040
rect 19616 32988 19668 33040
rect 12164 32852 12216 32904
rect 13636 32852 13688 32904
rect 16580 32852 16632 32904
rect 6552 32784 6604 32836
rect 8668 32784 8720 32836
rect 16212 32784 16264 32836
rect 20352 32963 20404 32972
rect 20352 32929 20361 32963
rect 20361 32929 20395 32963
rect 20395 32929 20404 32963
rect 20352 32920 20404 32929
rect 22468 32920 22520 32972
rect 23112 32920 23164 32972
rect 23388 32920 23440 32972
rect 19156 32852 19208 32904
rect 23296 32852 23348 32904
rect 24860 32852 24912 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 19064 32784 19116 32836
rect 6828 32716 6880 32768
rect 9312 32716 9364 32768
rect 12072 32716 12124 32768
rect 13268 32759 13320 32768
rect 13268 32725 13277 32759
rect 13277 32725 13311 32759
rect 13311 32725 13320 32759
rect 13268 32716 13320 32725
rect 14740 32716 14792 32768
rect 17040 32716 17092 32768
rect 20720 32784 20772 32836
rect 21916 32784 21968 32836
rect 23020 32827 23072 32836
rect 23020 32793 23029 32827
rect 23029 32793 23063 32827
rect 23063 32793 23072 32827
rect 23020 32784 23072 32793
rect 21548 32716 21600 32768
rect 22560 32759 22612 32768
rect 22560 32725 22569 32759
rect 22569 32725 22603 32759
rect 22603 32725 22612 32759
rect 22560 32716 22612 32725
rect 23572 32716 23624 32768
rect 25136 32759 25188 32768
rect 25136 32725 25145 32759
rect 25145 32725 25179 32759
rect 25179 32725 25188 32759
rect 25136 32716 25188 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 8576 32512 8628 32564
rect 9496 32444 9548 32496
rect 940 32376 992 32428
rect 7748 32376 7800 32428
rect 10508 32376 10560 32428
rect 8668 32351 8720 32360
rect 8668 32317 8677 32351
rect 8677 32317 8711 32351
rect 8711 32317 8720 32351
rect 8668 32308 8720 32317
rect 1584 32215 1636 32224
rect 1584 32181 1593 32215
rect 1593 32181 1627 32215
rect 1627 32181 1636 32215
rect 1584 32172 1636 32181
rect 7656 32215 7708 32224
rect 7656 32181 7665 32215
rect 7665 32181 7699 32215
rect 7699 32181 7708 32215
rect 7656 32172 7708 32181
rect 9772 32172 9824 32224
rect 14832 32512 14884 32564
rect 17316 32555 17368 32564
rect 17316 32521 17325 32555
rect 17325 32521 17359 32555
rect 17359 32521 17368 32555
rect 17316 32512 17368 32521
rect 19340 32512 19392 32564
rect 19708 32512 19760 32564
rect 21272 32512 21324 32564
rect 22284 32512 22336 32564
rect 25136 32512 25188 32564
rect 16764 32444 16816 32496
rect 17408 32444 17460 32496
rect 20812 32444 20864 32496
rect 21364 32444 21416 32496
rect 13268 32376 13320 32428
rect 15844 32376 15896 32428
rect 14464 32351 14516 32360
rect 14464 32317 14473 32351
rect 14473 32317 14507 32351
rect 14507 32317 14516 32351
rect 14464 32308 14516 32317
rect 16764 32308 16816 32360
rect 18420 32376 18472 32428
rect 20260 32376 20312 32428
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 23296 32376 23348 32428
rect 25412 32376 25464 32428
rect 18972 32308 19024 32360
rect 17040 32240 17092 32292
rect 17408 32240 17460 32292
rect 17592 32240 17644 32292
rect 20812 32308 20864 32360
rect 23204 32351 23256 32360
rect 23204 32317 23213 32351
rect 23213 32317 23247 32351
rect 23247 32317 23256 32351
rect 23204 32308 23256 32317
rect 20996 32240 21048 32292
rect 12348 32172 12400 32224
rect 14280 32172 14332 32224
rect 14556 32172 14608 32224
rect 16304 32172 16356 32224
rect 17776 32172 17828 32224
rect 18420 32172 18472 32224
rect 19340 32172 19392 32224
rect 20444 32172 20496 32224
rect 20536 32215 20588 32224
rect 20536 32181 20545 32215
rect 20545 32181 20579 32215
rect 20579 32181 20588 32215
rect 20536 32172 20588 32181
rect 22008 32215 22060 32224
rect 22008 32181 22017 32215
rect 22017 32181 22051 32215
rect 22051 32181 22060 32215
rect 22008 32172 22060 32181
rect 22192 32172 22244 32224
rect 22836 32172 22888 32224
rect 23480 32172 23532 32224
rect 24308 32172 24360 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 6920 32011 6972 32020
rect 6920 31977 6929 32011
rect 6929 31977 6963 32011
rect 6963 31977 6972 32011
rect 6920 31968 6972 31977
rect 7840 31968 7892 32020
rect 9404 31968 9456 32020
rect 11060 31968 11112 32020
rect 11980 31968 12032 32020
rect 4896 31832 4948 31884
rect 8392 31832 8444 31884
rect 8484 31832 8536 31884
rect 9496 31832 9548 31884
rect 4712 31807 4764 31816
rect 4712 31773 4721 31807
rect 4721 31773 4755 31807
rect 4755 31773 4764 31807
rect 4712 31764 4764 31773
rect 6552 31764 6604 31816
rect 8944 31764 8996 31816
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 10508 31764 10560 31816
rect 7840 31671 7892 31680
rect 7840 31637 7849 31671
rect 7849 31637 7883 31671
rect 7883 31637 7892 31671
rect 7840 31628 7892 31637
rect 10324 31628 10376 31680
rect 12716 31832 12768 31884
rect 19984 31968 20036 32020
rect 20352 31968 20404 32020
rect 21364 31968 21416 32020
rect 16488 31900 16540 31952
rect 14464 31832 14516 31884
rect 16856 31832 16908 31884
rect 17224 31900 17276 31952
rect 17500 31900 17552 31952
rect 17776 31875 17828 31884
rect 17776 31841 17785 31875
rect 17785 31841 17819 31875
rect 17819 31841 17828 31875
rect 17776 31832 17828 31841
rect 17868 31875 17920 31884
rect 17868 31841 17877 31875
rect 17877 31841 17911 31875
rect 17911 31841 17920 31875
rect 17868 31832 17920 31841
rect 20444 31900 20496 31952
rect 21732 31900 21784 31952
rect 22284 31900 22336 31952
rect 23296 31900 23348 31952
rect 24676 31900 24728 31952
rect 20996 31832 21048 31884
rect 21088 31832 21140 31884
rect 23020 31832 23072 31884
rect 23480 31832 23532 31884
rect 15292 31696 15344 31748
rect 15384 31739 15436 31748
rect 15384 31705 15393 31739
rect 15393 31705 15427 31739
rect 15427 31705 15436 31739
rect 15384 31696 15436 31705
rect 12716 31671 12768 31680
rect 12716 31637 12725 31671
rect 12725 31637 12759 31671
rect 12759 31637 12768 31671
rect 12716 31628 12768 31637
rect 15200 31628 15252 31680
rect 15844 31696 15896 31748
rect 18696 31696 18748 31748
rect 20628 31696 20680 31748
rect 21916 31764 21968 31816
rect 24032 31807 24084 31816
rect 24032 31773 24041 31807
rect 24041 31773 24075 31807
rect 24075 31773 24084 31807
rect 24032 31764 24084 31773
rect 21456 31696 21508 31748
rect 16764 31628 16816 31680
rect 19708 31628 19760 31680
rect 20076 31628 20128 31680
rect 25596 31696 25648 31748
rect 22928 31628 22980 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 4620 31424 4672 31476
rect 4712 31424 4764 31476
rect 7012 31467 7064 31476
rect 7012 31433 7021 31467
rect 7021 31433 7055 31467
rect 7055 31433 7064 31467
rect 7012 31424 7064 31433
rect 10048 31424 10100 31476
rect 10784 31424 10836 31476
rect 17132 31424 17184 31476
rect 5080 31356 5132 31408
rect 19432 31356 19484 31408
rect 4160 31288 4212 31340
rect 5356 31220 5408 31272
rect 7380 31331 7432 31340
rect 7380 31297 7389 31331
rect 7389 31297 7423 31331
rect 7423 31297 7432 31331
rect 7380 31288 7432 31297
rect 7840 31288 7892 31340
rect 7472 31263 7524 31272
rect 7472 31229 7481 31263
rect 7481 31229 7515 31263
rect 7515 31229 7524 31263
rect 7472 31220 7524 31229
rect 7564 31263 7616 31272
rect 7564 31229 7573 31263
rect 7573 31229 7607 31263
rect 7607 31229 7616 31263
rect 7564 31220 7616 31229
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 20812 31288 20864 31340
rect 25872 31356 25924 31408
rect 22836 31288 22888 31340
rect 24400 31288 24452 31340
rect 10692 31263 10744 31272
rect 10692 31229 10701 31263
rect 10701 31229 10735 31263
rect 10735 31229 10744 31263
rect 10692 31220 10744 31229
rect 15292 31220 15344 31272
rect 5448 31152 5500 31204
rect 10508 31152 10560 31204
rect 18788 31152 18840 31204
rect 21456 31152 21508 31204
rect 25228 31152 25280 31204
rect 23848 31084 23900 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 7380 30880 7432 30932
rect 11244 30880 11296 30932
rect 13360 30880 13412 30932
rect 7748 30812 7800 30864
rect 12256 30812 12308 30864
rect 6276 30744 6328 30796
rect 7196 30744 7248 30796
rect 7656 30676 7708 30728
rect 9128 30744 9180 30796
rect 10324 30608 10376 30660
rect 17040 30812 17092 30864
rect 17316 30744 17368 30796
rect 25964 30812 26016 30864
rect 22652 30744 22704 30796
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 17408 30719 17460 30728
rect 17408 30685 17417 30719
rect 17417 30685 17451 30719
rect 17451 30685 17460 30719
rect 17408 30676 17460 30685
rect 24216 30744 24268 30796
rect 24492 30744 24544 30796
rect 9404 30540 9456 30592
rect 14464 30608 14516 30660
rect 15200 30608 15252 30660
rect 22468 30608 22520 30660
rect 24492 30608 24544 30660
rect 12532 30583 12584 30592
rect 12532 30549 12541 30583
rect 12541 30549 12575 30583
rect 12575 30549 12584 30583
rect 12532 30540 12584 30549
rect 12624 30540 12676 30592
rect 13360 30583 13412 30592
rect 13360 30549 13369 30583
rect 13369 30549 13403 30583
rect 13403 30549 13412 30583
rect 13360 30540 13412 30549
rect 14188 30540 14240 30592
rect 15936 30540 15988 30592
rect 16212 30540 16264 30592
rect 16672 30540 16724 30592
rect 24032 30583 24084 30592
rect 24032 30549 24041 30583
rect 24041 30549 24075 30583
rect 24075 30549 24084 30583
rect 24032 30540 24084 30549
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 9036 30336 9088 30388
rect 13360 30336 13412 30388
rect 16948 30336 17000 30388
rect 25044 30336 25096 30388
rect 10324 30268 10376 30320
rect 15016 30268 15068 30320
rect 18512 30268 18564 30320
rect 18604 30268 18656 30320
rect 18972 30268 19024 30320
rect 19892 30268 19944 30320
rect 20444 30268 20496 30320
rect 20812 30311 20864 30320
rect 20812 30277 20821 30311
rect 20821 30277 20855 30311
rect 20855 30277 20864 30311
rect 20812 30268 20864 30277
rect 21364 30268 21416 30320
rect 22284 30268 22336 30320
rect 24216 30268 24268 30320
rect 12992 30243 13044 30252
rect 12992 30209 13001 30243
rect 13001 30209 13035 30243
rect 13035 30209 13044 30243
rect 12992 30200 13044 30209
rect 14372 30200 14424 30252
rect 19156 30200 19208 30252
rect 8024 30175 8076 30184
rect 8024 30141 8033 30175
rect 8033 30141 8067 30175
rect 8067 30141 8076 30175
rect 8024 30132 8076 30141
rect 8392 30132 8444 30184
rect 9680 30132 9732 30184
rect 10416 30064 10468 30116
rect 14648 30132 14700 30184
rect 15292 30175 15344 30184
rect 15292 30141 15301 30175
rect 15301 30141 15335 30175
rect 15335 30141 15344 30175
rect 15292 30132 15344 30141
rect 14004 30064 14056 30116
rect 16948 30132 17000 30184
rect 17592 30132 17644 30184
rect 20168 30200 20220 30252
rect 21732 30200 21784 30252
rect 3608 29996 3660 30048
rect 8484 29996 8536 30048
rect 9404 29996 9456 30048
rect 10968 29996 11020 30048
rect 13544 29996 13596 30048
rect 14924 29996 14976 30048
rect 17316 29996 17368 30048
rect 20260 30132 20312 30184
rect 18512 30064 18564 30116
rect 19432 30064 19484 30116
rect 22652 30200 22704 30252
rect 24032 30132 24084 30184
rect 22652 30064 22704 30116
rect 20444 30039 20496 30048
rect 20444 30005 20453 30039
rect 20453 30005 20487 30039
rect 20487 30005 20496 30039
rect 20444 29996 20496 30005
rect 23480 29996 23532 30048
rect 23756 29996 23808 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 8944 29792 8996 29844
rect 7564 29724 7616 29776
rect 9680 29724 9732 29776
rect 1308 29656 1360 29708
rect 8024 29656 8076 29708
rect 9772 29699 9824 29708
rect 9772 29665 9781 29699
rect 9781 29665 9815 29699
rect 9815 29665 9824 29699
rect 9772 29656 9824 29665
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 1860 29588 1912 29640
rect 9404 29588 9456 29640
rect 12624 29792 12676 29844
rect 13360 29792 13412 29844
rect 14096 29792 14148 29844
rect 14924 29792 14976 29844
rect 19248 29792 19300 29844
rect 10416 29724 10468 29776
rect 12164 29724 12216 29776
rect 10140 29656 10192 29708
rect 10600 29656 10652 29708
rect 11244 29699 11296 29708
rect 11244 29665 11253 29699
rect 11253 29665 11287 29699
rect 11287 29665 11296 29699
rect 11244 29656 11296 29665
rect 12440 29656 12492 29708
rect 13452 29699 13504 29708
rect 13452 29665 13461 29699
rect 13461 29665 13495 29699
rect 13495 29665 13504 29699
rect 13452 29656 13504 29665
rect 19616 29724 19668 29776
rect 20720 29724 20772 29776
rect 21272 29724 21324 29776
rect 3516 29520 3568 29572
rect 6000 29520 6052 29572
rect 8852 29520 8904 29572
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 10968 29588 11020 29597
rect 12164 29588 12216 29640
rect 12532 29520 12584 29572
rect 14832 29588 14884 29640
rect 19340 29656 19392 29708
rect 18696 29588 18748 29640
rect 21180 29699 21232 29708
rect 21180 29665 21189 29699
rect 21189 29665 21223 29699
rect 21223 29665 21232 29699
rect 21180 29656 21232 29665
rect 21732 29656 21784 29708
rect 22468 29792 22520 29844
rect 25136 29835 25188 29844
rect 25136 29801 25145 29835
rect 25145 29801 25179 29835
rect 25179 29801 25188 29835
rect 25136 29792 25188 29801
rect 24032 29724 24084 29776
rect 23480 29656 23532 29708
rect 23756 29699 23808 29708
rect 23756 29665 23765 29699
rect 23765 29665 23799 29699
rect 23799 29665 23808 29699
rect 23756 29656 23808 29665
rect 22192 29588 22244 29640
rect 22376 29631 22428 29640
rect 22376 29597 22385 29631
rect 22385 29597 22419 29631
rect 22419 29597 22428 29631
rect 22376 29588 22428 29597
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 12900 29452 12952 29504
rect 18328 29520 18380 29572
rect 23572 29520 23624 29572
rect 17500 29495 17552 29504
rect 17500 29461 17509 29495
rect 17509 29461 17543 29495
rect 17543 29461 17552 29495
rect 17500 29452 17552 29461
rect 17592 29495 17644 29504
rect 17592 29461 17601 29495
rect 17601 29461 17635 29495
rect 17635 29461 17644 29495
rect 17592 29452 17644 29461
rect 18972 29452 19024 29504
rect 19340 29452 19392 29504
rect 19984 29452 20036 29504
rect 20996 29452 21048 29504
rect 23296 29452 23348 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8208 29248 8260 29300
rect 12440 29248 12492 29300
rect 13360 29248 13412 29300
rect 13728 29248 13780 29300
rect 17500 29248 17552 29300
rect 8668 29180 8720 29232
rect 10324 29180 10376 29232
rect 11152 29180 11204 29232
rect 14372 29180 14424 29232
rect 17132 29180 17184 29232
rect 14556 29155 14608 29164
rect 14556 29121 14565 29155
rect 14565 29121 14599 29155
rect 14599 29121 14608 29155
rect 14556 29112 14608 29121
rect 19064 29180 19116 29232
rect 19524 29248 19576 29300
rect 21088 29248 21140 29300
rect 20628 29180 20680 29232
rect 24584 29180 24636 29232
rect 9680 29044 9732 29096
rect 10232 28976 10284 29028
rect 12440 28976 12492 29028
rect 12624 28976 12676 29028
rect 12900 28976 12952 29028
rect 14924 28976 14976 29028
rect 15844 29019 15896 29028
rect 15844 28985 15853 29019
rect 15853 28985 15887 29019
rect 15887 28985 15896 29019
rect 15844 28976 15896 28985
rect 16028 28976 16080 29028
rect 16764 28976 16816 29028
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 18144 29044 18196 29096
rect 19064 28976 19116 29028
rect 24400 28976 24452 29028
rect 11060 28908 11112 28960
rect 18604 28908 18656 28960
rect 22192 28951 22244 28960
rect 22192 28917 22201 28951
rect 22201 28917 22235 28951
rect 22235 28917 22244 28951
rect 22192 28908 22244 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 9312 28704 9364 28756
rect 9588 28704 9640 28756
rect 15384 28704 15436 28756
rect 16304 28747 16356 28756
rect 16304 28713 16313 28747
rect 16313 28713 16347 28747
rect 16347 28713 16356 28747
rect 16304 28704 16356 28713
rect 16488 28704 16540 28756
rect 20812 28704 20864 28756
rect 23296 28704 23348 28756
rect 23940 28704 23992 28756
rect 3424 28568 3476 28620
rect 6920 28568 6972 28620
rect 8208 28568 8260 28620
rect 8576 28568 8628 28620
rect 16396 28636 16448 28688
rect 12532 28568 12584 28620
rect 14280 28568 14332 28620
rect 17868 28568 17920 28620
rect 20720 28568 20772 28620
rect 20904 28568 20956 28620
rect 21180 28611 21232 28620
rect 21180 28577 21189 28611
rect 21189 28577 21223 28611
rect 21223 28577 21232 28611
rect 21180 28568 21232 28577
rect 22652 28568 22704 28620
rect 6276 28543 6328 28552
rect 6276 28509 6285 28543
rect 6285 28509 6319 28543
rect 6319 28509 6328 28543
rect 6276 28500 6328 28509
rect 8668 28500 8720 28552
rect 11244 28543 11296 28552
rect 11244 28509 11253 28543
rect 11253 28509 11287 28543
rect 11287 28509 11296 28543
rect 11244 28500 11296 28509
rect 12624 28500 12676 28552
rect 19984 28500 20036 28552
rect 20352 28500 20404 28552
rect 5816 28475 5868 28484
rect 5816 28441 5825 28475
rect 5825 28441 5859 28475
rect 5859 28441 5868 28475
rect 5816 28432 5868 28441
rect 7288 28432 7340 28484
rect 3976 28364 4028 28416
rect 4068 28364 4120 28416
rect 8760 28432 8812 28484
rect 15384 28432 15436 28484
rect 22192 28543 22244 28552
rect 22192 28509 22201 28543
rect 22201 28509 22235 28543
rect 22235 28509 22244 28543
rect 22192 28500 22244 28509
rect 24860 28500 24912 28552
rect 25320 28543 25372 28552
rect 25320 28509 25329 28543
rect 25329 28509 25363 28543
rect 25363 28509 25372 28543
rect 25320 28500 25372 28509
rect 8300 28364 8352 28416
rect 12808 28364 12860 28416
rect 16948 28407 17000 28416
rect 16948 28373 16957 28407
rect 16957 28373 16991 28407
rect 16991 28373 17000 28407
rect 16948 28364 17000 28373
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 20812 28364 20864 28416
rect 22652 28364 22704 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 7840 28160 7892 28212
rect 9680 28160 9732 28212
rect 10324 28160 10376 28212
rect 7288 28092 7340 28144
rect 8668 28024 8720 28076
rect 11060 28160 11112 28212
rect 12348 28203 12400 28212
rect 12348 28169 12357 28203
rect 12357 28169 12391 28203
rect 12391 28169 12400 28203
rect 12348 28160 12400 28169
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 17408 28160 17460 28212
rect 11888 28092 11940 28144
rect 13360 28092 13412 28144
rect 12624 28024 12676 28076
rect 14096 28024 14148 28076
rect 14280 28024 14332 28076
rect 18328 28024 18380 28076
rect 18880 28092 18932 28144
rect 20536 28092 20588 28144
rect 6276 27956 6328 28008
rect 8300 27956 8352 28008
rect 10784 27956 10836 28008
rect 10876 27888 10928 27940
rect 7564 27820 7616 27872
rect 12348 27820 12400 27872
rect 14372 27888 14424 27940
rect 16764 27956 16816 28008
rect 18420 27956 18472 28008
rect 18604 27999 18656 28008
rect 18604 27965 18613 27999
rect 18613 27965 18647 27999
rect 18647 27965 18656 27999
rect 18604 27956 18656 27965
rect 15108 27888 15160 27940
rect 19432 28024 19484 28076
rect 22560 28160 22612 28212
rect 23664 28092 23716 28144
rect 19248 27956 19300 28008
rect 20076 27999 20128 28008
rect 20076 27965 20085 27999
rect 20085 27965 20119 27999
rect 20119 27965 20128 27999
rect 20076 27956 20128 27965
rect 22836 28024 22888 28076
rect 23480 28067 23532 28076
rect 23480 28033 23489 28067
rect 23489 28033 23523 28067
rect 23523 28033 23532 28067
rect 23480 28024 23532 28033
rect 24032 28024 24084 28076
rect 23756 27956 23808 28008
rect 22100 27888 22152 27940
rect 13360 27863 13412 27872
rect 13360 27829 13369 27863
rect 13369 27829 13403 27863
rect 13403 27829 13412 27863
rect 13360 27820 13412 27829
rect 16580 27820 16632 27872
rect 19892 27820 19944 27872
rect 21916 27820 21968 27872
rect 23296 27863 23348 27872
rect 23296 27829 23305 27863
rect 23305 27829 23339 27863
rect 23339 27829 23348 27863
rect 23296 27820 23348 27829
rect 23940 27863 23992 27872
rect 23940 27829 23949 27863
rect 23949 27829 23983 27863
rect 23983 27829 23992 27863
rect 23940 27820 23992 27829
rect 24216 27820 24268 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 7840 27616 7892 27668
rect 12624 27616 12676 27668
rect 13084 27616 13136 27668
rect 15292 27616 15344 27668
rect 23296 27616 23348 27668
rect 12532 27548 12584 27600
rect 1308 27480 1360 27532
rect 3332 27480 3384 27532
rect 14464 27480 14516 27532
rect 14740 27523 14792 27532
rect 14740 27489 14749 27523
rect 14749 27489 14783 27523
rect 14783 27489 14792 27523
rect 14740 27480 14792 27489
rect 15936 27480 15988 27532
rect 16304 27548 16356 27600
rect 17040 27480 17092 27532
rect 17224 27523 17276 27532
rect 17224 27489 17233 27523
rect 17233 27489 17267 27523
rect 17267 27489 17276 27523
rect 17224 27480 17276 27489
rect 19524 27548 19576 27600
rect 23756 27548 23808 27600
rect 18420 27523 18472 27532
rect 18420 27489 18429 27523
rect 18429 27489 18463 27523
rect 18463 27489 18472 27523
rect 18420 27480 18472 27489
rect 18512 27523 18564 27532
rect 18512 27489 18521 27523
rect 18521 27489 18555 27523
rect 18555 27489 18564 27523
rect 18512 27480 18564 27489
rect 23296 27480 23348 27532
rect 1952 27412 2004 27464
rect 6276 27455 6328 27464
rect 6276 27421 6285 27455
rect 6285 27421 6319 27455
rect 6319 27421 6328 27455
rect 6276 27412 6328 27421
rect 10508 27412 10560 27464
rect 13176 27412 13228 27464
rect 16948 27412 17000 27464
rect 17960 27412 18012 27464
rect 22192 27412 22244 27464
rect 23848 27412 23900 27464
rect 6092 27344 6144 27396
rect 7288 27344 7340 27396
rect 4068 27276 4120 27328
rect 8392 27276 8444 27328
rect 15660 27344 15712 27396
rect 16120 27344 16172 27396
rect 18604 27344 18656 27396
rect 22468 27344 22520 27396
rect 24124 27344 24176 27396
rect 24860 27387 24912 27396
rect 24860 27353 24869 27387
rect 24869 27353 24903 27387
rect 24903 27353 24912 27387
rect 24860 27344 24912 27353
rect 13176 27319 13228 27328
rect 13176 27285 13185 27319
rect 13185 27285 13219 27319
rect 13219 27285 13228 27319
rect 13176 27276 13228 27285
rect 13912 27276 13964 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 16028 27319 16080 27328
rect 16028 27285 16037 27319
rect 16037 27285 16071 27319
rect 16071 27285 16080 27319
rect 16028 27276 16080 27285
rect 17224 27276 17276 27328
rect 17776 27276 17828 27328
rect 23848 27276 23900 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 1768 27072 1820 27124
rect 3516 27072 3568 27124
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 10784 27072 10836 27124
rect 14004 27072 14056 27124
rect 15108 27072 15160 27124
rect 15752 27072 15804 27124
rect 5908 27004 5960 27056
rect 6092 27004 6144 27056
rect 12072 27004 12124 27056
rect 2872 26936 2924 26988
rect 3608 26936 3660 26988
rect 9312 26936 9364 26988
rect 9404 26936 9456 26988
rect 11244 26936 11296 26988
rect 11428 26936 11480 26988
rect 13084 26936 13136 26988
rect 14004 26936 14056 26988
rect 14096 26936 14148 26988
rect 17500 27072 17552 27124
rect 17868 27115 17920 27124
rect 17868 27081 17877 27115
rect 17877 27081 17911 27115
rect 17911 27081 17920 27115
rect 17868 27072 17920 27081
rect 16028 27004 16080 27056
rect 18788 27004 18840 27056
rect 20352 27072 20404 27124
rect 22192 27072 22244 27124
rect 22468 27072 22520 27124
rect 19616 27047 19668 27056
rect 19616 27013 19625 27047
rect 19625 27013 19659 27047
rect 19659 27013 19668 27047
rect 19616 27004 19668 27013
rect 21272 27004 21324 27056
rect 24124 27004 24176 27056
rect 24676 27047 24728 27056
rect 24676 27013 24685 27047
rect 24685 27013 24719 27047
rect 24719 27013 24728 27047
rect 24676 27004 24728 27013
rect 7380 26868 7432 26920
rect 4896 26732 4948 26784
rect 7748 26800 7800 26852
rect 7840 26800 7892 26852
rect 8300 26868 8352 26920
rect 13452 26868 13504 26920
rect 15108 26911 15160 26920
rect 15108 26877 15117 26911
rect 15117 26877 15151 26911
rect 15151 26877 15160 26911
rect 15108 26868 15160 26877
rect 12992 26800 13044 26852
rect 17132 26800 17184 26852
rect 18696 26868 18748 26920
rect 19708 26868 19760 26920
rect 20076 26868 20128 26920
rect 20628 26868 20680 26920
rect 22192 26911 22244 26920
rect 22192 26877 22201 26911
rect 22201 26877 22235 26911
rect 22235 26877 22244 26911
rect 22192 26868 22244 26877
rect 22468 26911 22520 26920
rect 22468 26877 22477 26911
rect 22477 26877 22511 26911
rect 22511 26877 22520 26911
rect 22468 26868 22520 26877
rect 7012 26732 7064 26784
rect 7288 26732 7340 26784
rect 8576 26732 8628 26784
rect 8944 26775 8996 26784
rect 8944 26741 8953 26775
rect 8953 26741 8987 26775
rect 8987 26741 8996 26775
rect 8944 26732 8996 26741
rect 11980 26732 12032 26784
rect 14648 26775 14700 26784
rect 14648 26741 14657 26775
rect 14657 26741 14691 26775
rect 14691 26741 14700 26775
rect 14648 26732 14700 26741
rect 17408 26775 17460 26784
rect 17408 26741 17417 26775
rect 17417 26741 17451 26775
rect 17451 26741 17460 26775
rect 17408 26732 17460 26741
rect 20260 26732 20312 26784
rect 23204 26732 23256 26784
rect 23572 26732 23624 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 7104 26528 7156 26580
rect 7564 26528 7616 26580
rect 9312 26571 9364 26580
rect 9312 26537 9321 26571
rect 9321 26537 9355 26571
rect 9355 26537 9364 26571
rect 9312 26528 9364 26537
rect 11060 26528 11112 26580
rect 7748 26460 7800 26512
rect 10048 26460 10100 26512
rect 1584 26392 1636 26444
rect 4896 26435 4948 26444
rect 4896 26401 4905 26435
rect 4905 26401 4939 26435
rect 4939 26401 4948 26435
rect 4896 26392 4948 26401
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 10784 26435 10836 26444
rect 10784 26401 10793 26435
rect 10793 26401 10827 26435
rect 10827 26401 10836 26435
rect 10784 26392 10836 26401
rect 8392 26324 8444 26376
rect 10508 26367 10560 26376
rect 10508 26333 10517 26367
rect 10517 26333 10551 26367
rect 10551 26333 10560 26367
rect 10508 26324 10560 26333
rect 13176 26528 13228 26580
rect 14004 26528 14056 26580
rect 15384 26528 15436 26580
rect 16028 26528 16080 26580
rect 16212 26571 16264 26580
rect 16212 26537 16221 26571
rect 16221 26537 16255 26571
rect 16255 26537 16264 26571
rect 16212 26528 16264 26537
rect 16764 26528 16816 26580
rect 22376 26528 22428 26580
rect 23296 26528 23348 26580
rect 23848 26571 23900 26580
rect 23848 26537 23857 26571
rect 23857 26537 23891 26571
rect 23891 26537 23900 26571
rect 23848 26528 23900 26537
rect 13728 26460 13780 26512
rect 14188 26392 14240 26444
rect 17776 26392 17828 26444
rect 20260 26392 20312 26444
rect 22192 26392 22244 26444
rect 22744 26392 22796 26444
rect 13544 26324 13596 26376
rect 14464 26367 14516 26376
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 24952 26324 25004 26376
rect 3884 26256 3936 26308
rect 6460 26256 6512 26308
rect 7288 26256 7340 26308
rect 10600 26299 10652 26308
rect 10600 26265 10609 26299
rect 10609 26265 10643 26299
rect 10643 26265 10652 26299
rect 10600 26256 10652 26265
rect 16028 26256 16080 26308
rect 16856 26256 16908 26308
rect 19984 26256 20036 26308
rect 21640 26256 21692 26308
rect 16396 26188 16448 26240
rect 16764 26188 16816 26240
rect 17316 26188 17368 26240
rect 21272 26188 21324 26240
rect 24124 26256 24176 26308
rect 24308 26256 24360 26308
rect 25044 26256 25096 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 3976 25984 4028 26036
rect 8944 25984 8996 26036
rect 10232 25984 10284 26036
rect 15292 25984 15344 26036
rect 19432 25984 19484 26036
rect 19524 26027 19576 26036
rect 19524 25993 19533 26027
rect 19533 25993 19567 26027
rect 19567 25993 19576 26027
rect 19524 25984 19576 25993
rect 21088 25984 21140 26036
rect 22008 25984 22060 26036
rect 22284 25984 22336 26036
rect 8576 25916 8628 25968
rect 15108 25959 15160 25968
rect 15108 25925 15117 25959
rect 15117 25925 15151 25959
rect 15151 25925 15160 25959
rect 15108 25916 15160 25925
rect 16764 25916 16816 25968
rect 17868 25916 17920 25968
rect 25228 25916 25280 25968
rect 3332 25848 3384 25900
rect 3424 25848 3476 25900
rect 6920 25848 6972 25900
rect 3608 25780 3660 25832
rect 2872 25712 2924 25764
rect 3792 25712 3844 25764
rect 7196 25780 7248 25832
rect 13176 25848 13228 25900
rect 20444 25848 20496 25900
rect 22284 25848 22336 25900
rect 8392 25780 8444 25832
rect 11428 25780 11480 25832
rect 11796 25823 11848 25832
rect 11796 25789 11805 25823
rect 11805 25789 11839 25823
rect 11839 25789 11848 25823
rect 11796 25780 11848 25789
rect 12808 25780 12860 25832
rect 16396 25780 16448 25832
rect 17776 25780 17828 25832
rect 19616 25780 19668 25832
rect 19708 25823 19760 25832
rect 19708 25789 19717 25823
rect 19717 25789 19751 25823
rect 19751 25789 19760 25823
rect 19708 25780 19760 25789
rect 21732 25780 21784 25832
rect 9404 25712 9456 25764
rect 7196 25644 7248 25696
rect 10600 25712 10652 25764
rect 13544 25687 13596 25696
rect 13544 25653 13553 25687
rect 13553 25653 13587 25687
rect 13587 25653 13596 25687
rect 13544 25644 13596 25653
rect 14556 25712 14608 25764
rect 21456 25712 21508 25764
rect 14924 25644 14976 25696
rect 15752 25644 15804 25696
rect 18696 25644 18748 25696
rect 19524 25644 19576 25696
rect 21732 25644 21784 25696
rect 22100 25644 22152 25696
rect 23296 25780 23348 25832
rect 23480 25712 23532 25764
rect 25228 25712 25280 25764
rect 22744 25644 22796 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 4620 25440 4672 25492
rect 5816 25440 5868 25492
rect 6276 25440 6328 25492
rect 15108 25440 15160 25492
rect 19616 25440 19668 25492
rect 19800 25440 19852 25492
rect 14556 25372 14608 25424
rect 1308 25304 1360 25356
rect 6460 25347 6512 25356
rect 6460 25313 6469 25347
rect 6469 25313 6503 25347
rect 6503 25313 6512 25347
rect 6460 25304 6512 25313
rect 7104 25304 7156 25356
rect 7472 25304 7524 25356
rect 12808 25347 12860 25356
rect 12808 25313 12817 25347
rect 12817 25313 12851 25347
rect 12851 25313 12860 25347
rect 12808 25304 12860 25313
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 15660 25347 15712 25356
rect 15660 25313 15669 25347
rect 15669 25313 15703 25347
rect 15703 25313 15712 25347
rect 15660 25304 15712 25313
rect 18328 25304 18380 25356
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 3700 25236 3752 25288
rect 3976 25279 4028 25288
rect 3976 25245 3985 25279
rect 3985 25245 4019 25279
rect 4019 25245 4028 25279
rect 3976 25236 4028 25245
rect 7840 25236 7892 25288
rect 9036 25236 9088 25288
rect 11336 25236 11388 25288
rect 14464 25236 14516 25288
rect 16856 25279 16908 25288
rect 16856 25245 16865 25279
rect 16865 25245 16899 25279
rect 16899 25245 16908 25279
rect 16856 25236 16908 25245
rect 20352 25347 20404 25356
rect 20352 25313 20361 25347
rect 20361 25313 20395 25347
rect 20395 25313 20404 25347
rect 20352 25304 20404 25313
rect 20628 25347 20680 25356
rect 20628 25313 20637 25347
rect 20637 25313 20671 25347
rect 20671 25313 20680 25347
rect 20628 25304 20680 25313
rect 22652 25304 22704 25356
rect 23388 25304 23440 25356
rect 23940 25236 23992 25288
rect 3608 25100 3660 25152
rect 8208 25143 8260 25152
rect 8208 25109 8217 25143
rect 8217 25109 8251 25143
rect 8251 25109 8260 25143
rect 8208 25100 8260 25109
rect 9772 25100 9824 25152
rect 11704 25100 11756 25152
rect 16304 25168 16356 25220
rect 19064 25168 19116 25220
rect 21272 25168 21324 25220
rect 22284 25168 22336 25220
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 16672 25100 16724 25152
rect 20812 25100 20864 25152
rect 20904 25100 20956 25152
rect 21640 25100 21692 25152
rect 22560 25143 22612 25152
rect 22560 25109 22569 25143
rect 22569 25109 22603 25143
rect 22603 25109 22612 25143
rect 22560 25100 22612 25109
rect 22652 25100 22704 25152
rect 24124 25100 24176 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 6000 24828 6052 24880
rect 6184 24828 6236 24880
rect 2872 24760 2924 24812
rect 7012 24896 7064 24948
rect 7840 24896 7892 24948
rect 10876 24939 10928 24948
rect 10876 24905 10885 24939
rect 10885 24905 10919 24939
rect 10919 24905 10928 24939
rect 10876 24896 10928 24905
rect 9496 24828 9548 24880
rect 9680 24760 9732 24812
rect 9864 24760 9916 24812
rect 12072 24939 12124 24948
rect 12072 24905 12081 24939
rect 12081 24905 12115 24939
rect 12115 24905 12124 24939
rect 12072 24896 12124 24905
rect 12440 24896 12492 24948
rect 13636 24896 13688 24948
rect 19340 24896 19392 24948
rect 19524 24939 19576 24948
rect 19524 24905 19533 24939
rect 19533 24905 19567 24939
rect 19567 24905 19576 24939
rect 19524 24896 19576 24905
rect 12532 24760 12584 24812
rect 12900 24760 12952 24812
rect 13360 24760 13412 24812
rect 13636 24760 13688 24812
rect 14464 24760 14516 24812
rect 15936 24760 15988 24812
rect 19432 24760 19484 24812
rect 22468 24896 22520 24948
rect 24032 24828 24084 24880
rect 2780 24692 2832 24744
rect 6000 24692 6052 24744
rect 6460 24692 6512 24744
rect 7012 24692 7064 24744
rect 8208 24735 8260 24744
rect 8208 24701 8217 24735
rect 8217 24701 8251 24735
rect 8251 24701 8260 24735
rect 8208 24692 8260 24701
rect 11060 24692 11112 24744
rect 16212 24692 16264 24744
rect 16304 24735 16356 24744
rect 16304 24701 16313 24735
rect 16313 24701 16347 24735
rect 16347 24701 16356 24735
rect 16304 24692 16356 24701
rect 17408 24692 17460 24744
rect 18604 24735 18656 24744
rect 18604 24701 18613 24735
rect 18613 24701 18647 24735
rect 18647 24701 18656 24735
rect 18604 24692 18656 24701
rect 20628 24692 20680 24744
rect 1952 24624 2004 24676
rect 9404 24624 9456 24676
rect 14372 24624 14424 24676
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 22376 24692 22428 24744
rect 22836 24692 22888 24744
rect 23664 24692 23716 24744
rect 3976 24556 4028 24608
rect 4436 24556 4488 24608
rect 4620 24556 4672 24608
rect 8208 24556 8260 24608
rect 15016 24556 15068 24608
rect 18420 24556 18472 24608
rect 19800 24556 19852 24608
rect 22100 24599 22152 24608
rect 22100 24565 22109 24599
rect 22109 24565 22143 24599
rect 22143 24565 22152 24599
rect 22100 24556 22152 24565
rect 22376 24556 22428 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 4068 24352 4120 24404
rect 9496 24352 9548 24404
rect 19432 24352 19484 24404
rect 22468 24352 22520 24404
rect 4252 24284 4304 24336
rect 13544 24284 13596 24336
rect 4436 24216 4488 24268
rect 7472 24216 7524 24268
rect 9404 24259 9456 24268
rect 9404 24225 9413 24259
rect 9413 24225 9447 24259
rect 9447 24225 9456 24259
rect 9404 24216 9456 24225
rect 12164 24259 12216 24268
rect 12164 24225 12173 24259
rect 12173 24225 12207 24259
rect 12207 24225 12216 24259
rect 12164 24216 12216 24225
rect 2228 24080 2280 24132
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 13452 24148 13504 24200
rect 14648 24216 14700 24268
rect 15752 24216 15804 24268
rect 16212 24216 16264 24268
rect 17684 24216 17736 24268
rect 18512 24216 18564 24268
rect 19892 24259 19944 24268
rect 19892 24225 19901 24259
rect 19901 24225 19935 24259
rect 19935 24225 19944 24259
rect 19892 24216 19944 24225
rect 20904 24216 20956 24268
rect 21088 24259 21140 24268
rect 21088 24225 21097 24259
rect 21097 24225 21131 24259
rect 21131 24225 21140 24259
rect 21088 24216 21140 24225
rect 21272 24259 21324 24268
rect 21272 24225 21281 24259
rect 21281 24225 21315 24259
rect 21315 24225 21324 24259
rect 21272 24216 21324 24225
rect 16672 24148 16724 24200
rect 19800 24191 19852 24200
rect 19800 24157 19809 24191
rect 19809 24157 19843 24191
rect 19843 24157 19852 24191
rect 19800 24148 19852 24157
rect 24400 24148 24452 24200
rect 24768 24148 24820 24200
rect 8484 24080 8536 24132
rect 9496 24080 9548 24132
rect 10416 24080 10468 24132
rect 13084 24080 13136 24132
rect 18880 24080 18932 24132
rect 24952 24080 25004 24132
rect 3424 24012 3476 24064
rect 8392 24012 8444 24064
rect 8760 24012 8812 24064
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 11520 24055 11572 24064
rect 11520 24021 11529 24055
rect 11529 24021 11563 24055
rect 11563 24021 11572 24055
rect 11520 24012 11572 24021
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 14556 24012 14608 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 17776 24055 17828 24064
rect 17776 24021 17785 24055
rect 17785 24021 17819 24055
rect 17819 24021 17828 24055
rect 17776 24012 17828 24021
rect 17868 24012 17920 24064
rect 18788 24012 18840 24064
rect 20628 24055 20680 24064
rect 20628 24021 20637 24055
rect 20637 24021 20671 24055
rect 20671 24021 20680 24055
rect 20628 24012 20680 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 2688 23808 2740 23860
rect 4068 23808 4120 23860
rect 5540 23808 5592 23860
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 9036 23808 9088 23860
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 13084 23851 13136 23860
rect 13084 23817 13093 23851
rect 13093 23817 13127 23851
rect 13127 23817 13136 23851
rect 13084 23808 13136 23817
rect 13452 23851 13504 23860
rect 13452 23817 13461 23851
rect 13461 23817 13495 23851
rect 13495 23817 13504 23851
rect 13452 23808 13504 23817
rect 13636 23808 13688 23860
rect 14188 23808 14240 23860
rect 21088 23808 21140 23860
rect 23480 23808 23532 23860
rect 4988 23740 5040 23792
rect 6644 23740 6696 23792
rect 11612 23740 11664 23792
rect 11980 23740 12032 23792
rect 4068 23672 4120 23724
rect 4620 23604 4672 23656
rect 4988 23604 5040 23656
rect 7104 23672 7156 23724
rect 9036 23647 9088 23656
rect 9036 23613 9045 23647
rect 9045 23613 9079 23647
rect 9079 23613 9088 23647
rect 9036 23604 9088 23613
rect 4252 23468 4304 23520
rect 5816 23468 5868 23520
rect 8484 23511 8536 23520
rect 8484 23477 8493 23511
rect 8493 23477 8527 23511
rect 8527 23477 8536 23511
rect 8484 23468 8536 23477
rect 13544 23672 13596 23724
rect 16488 23672 16540 23724
rect 24860 23740 24912 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 24124 23715 24176 23724
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 9496 23604 9548 23656
rect 9404 23536 9456 23588
rect 10876 23604 10928 23656
rect 16396 23604 16448 23656
rect 23388 23604 23440 23656
rect 11980 23536 12032 23588
rect 15292 23468 15344 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 3332 23264 3384 23316
rect 5816 23264 5868 23316
rect 6828 23264 6880 23316
rect 16212 23196 16264 23248
rect 1308 23128 1360 23180
rect 5540 23171 5592 23180
rect 5540 23137 5549 23171
rect 5549 23137 5583 23171
rect 5583 23137 5592 23171
rect 5540 23128 5592 23137
rect 7012 23128 7064 23180
rect 7840 23128 7892 23180
rect 10140 23171 10192 23180
rect 10140 23137 10149 23171
rect 10149 23137 10183 23171
rect 10183 23137 10192 23171
rect 10140 23128 10192 23137
rect 16304 23171 16356 23180
rect 16304 23137 16313 23171
rect 16313 23137 16347 23171
rect 16347 23137 16356 23171
rect 16304 23128 16356 23137
rect 18880 23264 18932 23316
rect 19524 23264 19576 23316
rect 20720 23264 20772 23316
rect 22744 23196 22796 23248
rect 18512 23128 18564 23180
rect 18880 23128 18932 23180
rect 21916 23171 21968 23180
rect 21916 23137 21925 23171
rect 21925 23137 21959 23171
rect 21959 23137 21968 23171
rect 21916 23128 21968 23137
rect 22376 23128 22428 23180
rect 2688 23060 2740 23112
rect 15476 23060 15528 23112
rect 16580 23060 16632 23112
rect 5724 22992 5776 23044
rect 7104 22992 7156 23044
rect 9680 22992 9732 23044
rect 13728 22992 13780 23044
rect 22100 23060 22152 23112
rect 23572 23060 23624 23112
rect 26056 22992 26108 23044
rect 8300 22924 8352 22976
rect 9036 22924 9088 22976
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 11428 22924 11480 22976
rect 12256 22924 12308 22976
rect 14464 22924 14516 22976
rect 16764 22924 16816 22976
rect 17224 22924 17276 22976
rect 17316 22967 17368 22976
rect 17316 22933 17325 22967
rect 17325 22933 17359 22967
rect 17359 22933 17368 22967
rect 17316 22924 17368 22933
rect 19248 22924 19300 22976
rect 21180 22924 21232 22976
rect 22100 22924 22152 22976
rect 22652 22924 22704 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1768 22720 1820 22772
rect 2872 22720 2924 22772
rect 3884 22720 3936 22772
rect 10048 22720 10100 22772
rect 14464 22720 14516 22772
rect 14556 22720 14608 22772
rect 15660 22720 15712 22772
rect 16396 22720 16448 22772
rect 9680 22652 9732 22704
rect 12624 22652 12676 22704
rect 13636 22695 13688 22704
rect 13636 22661 13645 22695
rect 13645 22661 13679 22695
rect 13679 22661 13688 22695
rect 13636 22652 13688 22661
rect 15936 22652 15988 22704
rect 16488 22652 16540 22704
rect 18512 22720 18564 22772
rect 19064 22652 19116 22704
rect 19800 22652 19852 22704
rect 22376 22720 22428 22772
rect 23480 22720 23532 22772
rect 2872 22584 2924 22636
rect 3516 22584 3568 22636
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 7656 22584 7708 22636
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 3424 22516 3476 22568
rect 6000 22516 6052 22568
rect 7840 22516 7892 22568
rect 4804 22448 4856 22500
rect 4160 22380 4212 22432
rect 10876 22516 10928 22568
rect 11796 22516 11848 22568
rect 12900 22584 12952 22636
rect 9128 22380 9180 22432
rect 12072 22448 12124 22500
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 13360 22559 13412 22568
rect 13360 22525 13369 22559
rect 13369 22525 13403 22559
rect 13403 22525 13412 22559
rect 13360 22516 13412 22525
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 10600 22423 10652 22432
rect 10600 22389 10609 22423
rect 10609 22389 10643 22423
rect 10643 22389 10652 22423
rect 10600 22380 10652 22389
rect 10968 22380 11020 22432
rect 12164 22423 12216 22432
rect 12164 22389 12173 22423
rect 12173 22389 12207 22423
rect 12207 22389 12216 22423
rect 12164 22380 12216 22389
rect 16764 22516 16816 22568
rect 17592 22516 17644 22568
rect 18972 22516 19024 22568
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 21272 22516 21324 22568
rect 24032 22652 24084 22704
rect 22192 22584 22244 22636
rect 22652 22516 22704 22568
rect 22836 22516 22888 22568
rect 15936 22380 15988 22432
rect 17132 22423 17184 22432
rect 17132 22389 17162 22423
rect 17162 22389 17184 22423
rect 17132 22380 17184 22389
rect 17684 22380 17736 22432
rect 18880 22380 18932 22432
rect 19064 22380 19116 22432
rect 19800 22380 19852 22432
rect 20352 22380 20404 22432
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 2688 22219 2740 22228
rect 2688 22185 2697 22219
rect 2697 22185 2731 22219
rect 2731 22185 2740 22219
rect 2688 22176 2740 22185
rect 5632 22176 5684 22228
rect 7472 22176 7524 22228
rect 3608 22040 3660 22092
rect 6828 22108 6880 22160
rect 7564 22108 7616 22160
rect 8944 22176 8996 22228
rect 10232 22176 10284 22228
rect 7104 22040 7156 22092
rect 7380 22040 7432 22092
rect 7472 22040 7524 22092
rect 11612 22108 11664 22160
rect 11796 22040 11848 22092
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 7012 21972 7064 22024
rect 9496 21972 9548 22024
rect 14280 22151 14332 22160
rect 14280 22117 14289 22151
rect 14289 22117 14323 22151
rect 14323 22117 14332 22151
rect 14280 22108 14332 22117
rect 12624 21972 12676 22024
rect 13636 22040 13688 22092
rect 18972 22176 19024 22228
rect 19064 22176 19116 22228
rect 22928 22176 22980 22228
rect 17684 22108 17736 22160
rect 16948 22040 17000 22092
rect 17776 22040 17828 22092
rect 19708 22108 19760 22160
rect 20076 22108 20128 22160
rect 22652 22108 22704 22160
rect 19616 22040 19668 22092
rect 13912 21972 13964 22024
rect 15200 21972 15252 22024
rect 17224 21972 17276 22024
rect 24216 21972 24268 22024
rect 8484 21904 8536 21956
rect 10048 21904 10100 21956
rect 15844 21904 15896 21956
rect 16028 21904 16080 21956
rect 16488 21904 16540 21956
rect 20352 21904 20404 21956
rect 24952 21904 25004 21956
rect 1768 21836 1820 21888
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 7288 21879 7340 21888
rect 7288 21845 7297 21879
rect 7297 21845 7331 21879
rect 7331 21845 7340 21879
rect 7288 21836 7340 21845
rect 7748 21879 7800 21888
rect 7748 21845 7757 21879
rect 7757 21845 7791 21879
rect 7791 21845 7800 21879
rect 7748 21836 7800 21845
rect 9496 21836 9548 21888
rect 12348 21879 12400 21888
rect 12348 21845 12357 21879
rect 12357 21845 12391 21879
rect 12391 21845 12400 21879
rect 12348 21836 12400 21845
rect 12716 21836 12768 21888
rect 13268 21836 13320 21888
rect 14648 21836 14700 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 14832 21836 14884 21888
rect 16120 21836 16172 21888
rect 17868 21836 17920 21888
rect 19892 21836 19944 21888
rect 20168 21836 20220 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 2964 21632 3016 21684
rect 5724 21632 5776 21684
rect 7288 21632 7340 21684
rect 7656 21632 7708 21684
rect 10692 21632 10744 21684
rect 14740 21632 14792 21684
rect 15200 21632 15252 21684
rect 17500 21632 17552 21684
rect 19340 21632 19392 21684
rect 2780 21564 2832 21616
rect 3332 21564 3384 21616
rect 9128 21564 9180 21616
rect 13268 21564 13320 21616
rect 13912 21564 13964 21616
rect 15844 21564 15896 21616
rect 18328 21564 18380 21616
rect 18972 21607 19024 21616
rect 18972 21573 18981 21607
rect 18981 21573 19015 21607
rect 19015 21573 19024 21607
rect 18972 21564 19024 21573
rect 19892 21607 19944 21616
rect 19892 21573 19901 21607
rect 19901 21573 19935 21607
rect 19935 21573 19944 21607
rect 19892 21564 19944 21573
rect 20352 21564 20404 21616
rect 3792 21496 3844 21548
rect 4160 21496 4212 21548
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 10232 21496 10284 21548
rect 11704 21496 11756 21548
rect 12348 21496 12400 21548
rect 12900 21496 12952 21548
rect 13728 21496 13780 21548
rect 2228 21428 2280 21480
rect 7196 21471 7248 21480
rect 7196 21437 7205 21471
rect 7205 21437 7239 21471
rect 7239 21437 7248 21471
rect 7196 21428 7248 21437
rect 7564 21360 7616 21412
rect 10416 21471 10468 21480
rect 10416 21437 10425 21471
rect 10425 21437 10459 21471
rect 10459 21437 10468 21471
rect 10416 21428 10468 21437
rect 10968 21428 11020 21480
rect 11980 21428 12032 21480
rect 13452 21428 13504 21480
rect 2780 21292 2832 21344
rect 5724 21292 5776 21344
rect 6184 21292 6236 21344
rect 12072 21360 12124 21412
rect 14924 21496 14976 21548
rect 17316 21496 17368 21548
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 21364 21496 21416 21548
rect 22836 21564 22888 21616
rect 23756 21632 23808 21684
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 14464 21471 14516 21480
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 19524 21360 19576 21412
rect 9680 21292 9732 21344
rect 13820 21292 13872 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 22192 21428 22244 21480
rect 22928 21428 22980 21480
rect 21548 21292 21600 21344
rect 24584 21292 24636 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 21088 2924 21140
rect 6552 21088 6604 21140
rect 8116 21088 8168 21140
rect 11980 21088 12032 21140
rect 13728 21131 13780 21140
rect 13728 21097 13737 21131
rect 13737 21097 13771 21131
rect 13771 21097 13780 21131
rect 13728 21088 13780 21097
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 3976 20995 4028 21004
rect 3976 20961 3985 20995
rect 3985 20961 4019 20995
rect 4019 20961 4028 20995
rect 3976 20952 4028 20961
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 10324 20952 10376 21004
rect 12072 20952 12124 21004
rect 12624 21020 12676 21072
rect 16672 21088 16724 21140
rect 21548 21088 21600 21140
rect 22376 21131 22428 21140
rect 22376 21097 22385 21131
rect 22385 21097 22419 21131
rect 22419 21097 22428 21131
rect 22376 21088 22428 21097
rect 13360 20952 13412 21004
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 19340 21020 19392 21072
rect 20536 21020 20588 21072
rect 18972 20952 19024 21004
rect 23480 20995 23532 21004
rect 23480 20961 23489 20995
rect 23489 20961 23523 20995
rect 23523 20961 23532 20995
rect 23480 20952 23532 20961
rect 2872 20884 2924 20936
rect 3516 20884 3568 20936
rect 11520 20884 11572 20936
rect 14188 20884 14240 20936
rect 16948 20927 17000 20936
rect 16948 20893 16957 20927
rect 16957 20893 16991 20927
rect 16991 20893 17000 20927
rect 16948 20884 17000 20893
rect 17868 20884 17920 20936
rect 19432 20884 19484 20936
rect 22192 20884 22244 20936
rect 22376 20884 22428 20936
rect 22744 20884 22796 20936
rect 5632 20816 5684 20868
rect 7656 20816 7708 20868
rect 16488 20816 16540 20868
rect 17500 20816 17552 20868
rect 20628 20816 20680 20868
rect 5724 20791 5776 20800
rect 5724 20757 5733 20791
rect 5733 20757 5767 20791
rect 5767 20757 5776 20791
rect 5724 20748 5776 20757
rect 6184 20748 6236 20800
rect 6368 20748 6420 20800
rect 6460 20748 6512 20800
rect 8576 20748 8628 20800
rect 9220 20748 9272 20800
rect 10692 20748 10744 20800
rect 11612 20748 11664 20800
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 16580 20748 16632 20800
rect 20352 20748 20404 20800
rect 21364 20816 21416 20868
rect 22928 20791 22980 20800
rect 22928 20757 22937 20791
rect 22937 20757 22971 20791
rect 22971 20757 22980 20791
rect 22928 20748 22980 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 7748 20544 7800 20596
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 12164 20544 12216 20596
rect 13820 20544 13872 20596
rect 15108 20544 15160 20596
rect 16948 20544 17000 20596
rect 17408 20544 17460 20596
rect 22928 20544 22980 20596
rect 23480 20544 23532 20596
rect 6828 20476 6880 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 7104 20408 7156 20460
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 8024 20408 8076 20460
rect 17040 20408 17092 20460
rect 18972 20476 19024 20528
rect 20352 20476 20404 20528
rect 20812 20476 20864 20528
rect 22560 20476 22612 20528
rect 23756 20476 23808 20528
rect 22652 20408 22704 20460
rect 1308 20340 1360 20392
rect 7932 20383 7984 20392
rect 7932 20349 7941 20383
rect 7941 20349 7975 20383
rect 7975 20349 7984 20383
rect 7932 20340 7984 20349
rect 12072 20340 12124 20392
rect 12164 20383 12216 20392
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 8576 20272 8628 20324
rect 10140 20272 10192 20324
rect 11060 20272 11112 20324
rect 13452 20340 13504 20392
rect 14464 20340 14516 20392
rect 16028 20340 16080 20392
rect 18512 20340 18564 20392
rect 20628 20272 20680 20324
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 11244 20204 11296 20256
rect 14740 20204 14792 20256
rect 15844 20204 15896 20256
rect 18236 20204 18288 20256
rect 20720 20204 20772 20256
rect 21640 20272 21692 20324
rect 22836 20204 22888 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 7012 20000 7064 20052
rect 7196 19864 7248 19916
rect 9128 20043 9180 20052
rect 9128 20009 9137 20043
rect 9137 20009 9171 20043
rect 9171 20009 9180 20043
rect 9128 20000 9180 20009
rect 12348 20000 12400 20052
rect 12900 20000 12952 20052
rect 21916 20000 21968 20052
rect 3332 19796 3384 19848
rect 1860 19660 1912 19712
rect 5632 19728 5684 19780
rect 5448 19660 5500 19712
rect 11244 19864 11296 19916
rect 11336 19864 11388 19916
rect 11152 19796 11204 19848
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 18420 19907 18472 19916
rect 18420 19873 18429 19907
rect 18429 19873 18463 19907
rect 18463 19873 18472 19907
rect 18420 19864 18472 19873
rect 20720 19932 20772 19984
rect 22652 19932 22704 19984
rect 24952 19864 25004 19916
rect 13360 19796 13412 19848
rect 14924 19796 14976 19848
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 18328 19796 18380 19848
rect 25228 19796 25280 19848
rect 6184 19728 6236 19780
rect 6828 19728 6880 19780
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 10140 19660 10192 19712
rect 11152 19660 11204 19712
rect 11704 19660 11756 19712
rect 12256 19660 12308 19712
rect 18604 19728 18656 19780
rect 19248 19728 19300 19780
rect 21824 19728 21876 19780
rect 18236 19660 18288 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 4804 19499 4856 19508
rect 4804 19465 4813 19499
rect 4813 19465 4847 19499
rect 4847 19465 4856 19499
rect 4804 19456 4856 19465
rect 7472 19456 7524 19508
rect 9680 19456 9732 19508
rect 10232 19456 10284 19508
rect 7840 19388 7892 19440
rect 11060 19456 11112 19508
rect 11612 19456 11664 19508
rect 15936 19456 15988 19508
rect 11796 19388 11848 19440
rect 12072 19388 12124 19440
rect 7564 19320 7616 19372
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 11704 19320 11756 19372
rect 9404 19252 9456 19304
rect 10324 19252 10376 19304
rect 17040 19388 17092 19440
rect 17224 19431 17276 19440
rect 17224 19397 17233 19431
rect 17233 19397 17267 19431
rect 17267 19397 17276 19431
rect 17224 19388 17276 19397
rect 20996 19456 21048 19508
rect 22192 19388 22244 19440
rect 24860 19388 24912 19440
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 15292 19320 15344 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 21088 19320 21140 19372
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 25044 19320 25096 19372
rect 12624 19252 12676 19304
rect 24676 19295 24728 19304
rect 24676 19261 24685 19295
rect 24685 19261 24719 19295
rect 24719 19261 24728 19295
rect 24676 19252 24728 19261
rect 23480 19184 23532 19236
rect 5632 19116 5684 19168
rect 6184 19116 6236 19168
rect 11336 19116 11388 19168
rect 12900 19116 12952 19168
rect 14464 19116 14516 19168
rect 17040 19116 17092 19168
rect 18972 19116 19024 19168
rect 20260 19116 20312 19168
rect 20444 19116 20496 19168
rect 22100 19116 22152 19168
rect 22376 19116 22428 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 3792 18912 3844 18964
rect 7012 18912 7064 18964
rect 8576 18912 8628 18964
rect 10968 18912 11020 18964
rect 3424 18776 3476 18828
rect 7748 18776 7800 18828
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 11612 18776 11664 18828
rect 12808 18776 12860 18828
rect 20444 18844 20496 18896
rect 22192 18844 22244 18896
rect 13452 18776 13504 18828
rect 17132 18776 17184 18828
rect 19248 18776 19300 18828
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 21364 18776 21416 18828
rect 22560 18776 22612 18828
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 5448 18751 5500 18760
rect 5448 18717 5457 18751
rect 5457 18717 5491 18751
rect 5491 18717 5500 18751
rect 5448 18708 5500 18717
rect 12716 18708 12768 18760
rect 14188 18708 14240 18760
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 18512 18708 18564 18760
rect 21732 18708 21784 18760
rect 22008 18708 22060 18760
rect 24584 18708 24636 18760
rect 1768 18572 1820 18624
rect 6184 18640 6236 18692
rect 12348 18640 12400 18692
rect 13544 18640 13596 18692
rect 19064 18640 19116 18692
rect 7840 18572 7892 18624
rect 11244 18572 11296 18624
rect 12072 18572 12124 18624
rect 15936 18572 15988 18624
rect 16580 18572 16632 18624
rect 20168 18572 20220 18624
rect 23756 18640 23808 18692
rect 22652 18572 22704 18624
rect 23296 18572 23348 18624
rect 24216 18572 24268 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 6184 18300 6236 18352
rect 1860 18232 1912 18284
rect 1308 18164 1360 18216
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 10600 18368 10652 18420
rect 11060 18411 11112 18420
rect 11060 18377 11069 18411
rect 11069 18377 11103 18411
rect 11103 18377 11112 18411
rect 11060 18368 11112 18377
rect 11704 18368 11756 18420
rect 13544 18368 13596 18420
rect 9680 18300 9732 18352
rect 10876 18300 10928 18352
rect 12348 18300 12400 18352
rect 18328 18300 18380 18352
rect 13728 18232 13780 18284
rect 18972 18232 19024 18284
rect 20904 18368 20956 18420
rect 23296 18368 23348 18420
rect 22468 18300 22520 18352
rect 22744 18300 22796 18352
rect 23756 18300 23808 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 22192 18232 22244 18284
rect 22376 18232 22428 18284
rect 7840 18028 7892 18080
rect 11336 18164 11388 18216
rect 12624 18164 12676 18216
rect 14464 18164 14516 18216
rect 17408 18164 17460 18216
rect 12164 18096 12216 18148
rect 22008 18164 22060 18216
rect 10232 18028 10284 18080
rect 13544 18028 13596 18080
rect 16580 18028 16632 18080
rect 20076 18028 20128 18080
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 22468 18096 22520 18148
rect 22652 18096 22704 18148
rect 23388 18028 23440 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 4436 17824 4488 17876
rect 5448 17688 5500 17740
rect 6184 17620 6236 17672
rect 6920 17620 6972 17672
rect 11520 17824 11572 17876
rect 16672 17824 16724 17876
rect 18788 17824 18840 17876
rect 19340 17824 19392 17876
rect 18420 17756 18472 17808
rect 20260 17824 20312 17876
rect 11980 17688 12032 17740
rect 13544 17688 13596 17740
rect 15476 17688 15528 17740
rect 17408 17688 17460 17740
rect 18788 17688 18840 17740
rect 19248 17688 19300 17740
rect 20352 17688 20404 17740
rect 14280 17620 14332 17672
rect 17316 17620 17368 17672
rect 19156 17620 19208 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 22284 17620 22336 17672
rect 7288 17552 7340 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 10232 17552 10284 17604
rect 6552 17527 6604 17536
rect 6552 17493 6561 17527
rect 6561 17493 6595 17527
rect 6595 17493 6604 17527
rect 6552 17484 6604 17493
rect 9588 17527 9640 17536
rect 9588 17493 9597 17527
rect 9597 17493 9631 17527
rect 9631 17493 9640 17527
rect 9588 17484 9640 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 14648 17527 14700 17536
rect 14648 17493 14657 17527
rect 14657 17493 14691 17527
rect 14691 17493 14700 17527
rect 14648 17484 14700 17493
rect 15108 17484 15160 17536
rect 18696 17552 18748 17604
rect 20720 17552 20772 17604
rect 19708 17484 19760 17536
rect 19984 17484 20036 17536
rect 20536 17484 20588 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 4160 17280 4212 17332
rect 5172 17212 5224 17264
rect 7012 17144 7064 17196
rect 7288 17212 7340 17264
rect 6552 17076 6604 17128
rect 7840 17008 7892 17060
rect 9864 17008 9916 17060
rect 9312 16940 9364 16992
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 12072 17323 12124 17332
rect 12072 17289 12081 17323
rect 12081 17289 12115 17323
rect 12115 17289 12124 17323
rect 12072 17280 12124 17289
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 14648 17280 14700 17332
rect 11704 17144 11756 17196
rect 13912 17212 13964 17264
rect 14740 17255 14792 17264
rect 14740 17221 14749 17255
rect 14749 17221 14783 17255
rect 14783 17221 14792 17255
rect 14740 17212 14792 17221
rect 15384 17280 15436 17332
rect 18420 17280 18472 17332
rect 19248 17280 19300 17332
rect 19432 17280 19484 17332
rect 17316 17212 17368 17264
rect 18144 17212 18196 17264
rect 11060 17076 11112 17128
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 15108 17144 15160 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 20904 17280 20956 17332
rect 19984 17255 20036 17264
rect 19984 17221 19993 17255
rect 19993 17221 20027 17255
rect 20027 17221 20036 17255
rect 19984 17212 20036 17221
rect 20720 17212 20772 17264
rect 21364 17280 21416 17332
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 12716 17008 12768 17060
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 14280 17076 14332 17128
rect 14464 17076 14516 17128
rect 17132 17076 17184 17128
rect 18420 17076 18472 17128
rect 22836 17076 22888 17128
rect 23756 17212 23808 17264
rect 13912 16940 13964 16992
rect 17776 16940 17828 16992
rect 22100 16940 22152 16992
rect 22744 16940 22796 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 2872 16736 2924 16788
rect 9588 16736 9640 16788
rect 10232 16736 10284 16788
rect 6552 16600 6604 16652
rect 7656 16600 7708 16652
rect 5632 16575 5684 16584
rect 5632 16541 5641 16575
rect 5641 16541 5675 16575
rect 5675 16541 5684 16575
rect 5632 16532 5684 16541
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 10324 16600 10376 16652
rect 10784 16643 10836 16652
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11336 16736 11388 16788
rect 12624 16736 12676 16788
rect 6184 16464 6236 16516
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 6920 16396 6972 16448
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9128 16532 9180 16584
rect 10876 16532 10928 16584
rect 12256 16600 12308 16652
rect 15476 16600 15528 16652
rect 22836 16600 22888 16652
rect 11336 16532 11388 16584
rect 16212 16532 16264 16584
rect 18328 16532 18380 16584
rect 21640 16532 21692 16584
rect 11060 16464 11112 16516
rect 20904 16464 20956 16516
rect 21916 16507 21968 16516
rect 21916 16473 21925 16507
rect 21925 16473 21959 16507
rect 21959 16473 21968 16507
rect 21916 16464 21968 16473
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 10876 16396 10928 16448
rect 12532 16396 12584 16448
rect 13544 16396 13596 16448
rect 15660 16396 15712 16448
rect 18144 16396 18196 16448
rect 18328 16396 18380 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 7012 16235 7064 16244
rect 7012 16201 7021 16235
rect 7021 16201 7055 16235
rect 7055 16201 7064 16235
rect 7012 16192 7064 16201
rect 7472 16235 7524 16244
rect 7472 16201 7481 16235
rect 7481 16201 7515 16235
rect 7515 16201 7524 16235
rect 7472 16192 7524 16201
rect 8576 16192 8628 16244
rect 9772 16192 9824 16244
rect 10876 16192 10928 16244
rect 18420 16192 18472 16244
rect 20444 16235 20496 16244
rect 20444 16201 20453 16235
rect 20453 16201 20487 16235
rect 20487 16201 20496 16235
rect 20444 16192 20496 16201
rect 23848 16192 23900 16244
rect 10692 16124 10744 16176
rect 14004 16124 14056 16176
rect 16120 16167 16172 16176
rect 16120 16133 16129 16167
rect 16129 16133 16163 16167
rect 16163 16133 16172 16167
rect 16120 16124 16172 16133
rect 17408 16124 17460 16176
rect 20996 16124 21048 16176
rect 22560 16124 22612 16176
rect 22744 16124 22796 16176
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 1308 15988 1360 16040
rect 7288 15988 7340 16040
rect 7656 15988 7708 16040
rect 12808 16056 12860 16108
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 10324 15988 10376 16040
rect 12348 15920 12400 15972
rect 7840 15852 7892 15904
rect 14832 15895 14884 15904
rect 14832 15861 14841 15895
rect 14841 15861 14875 15895
rect 14875 15861 14884 15895
rect 14832 15852 14884 15861
rect 15384 16056 15436 16108
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 20812 16056 20864 16108
rect 18328 15988 18380 16040
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 20904 15988 20956 16040
rect 16304 15963 16356 15972
rect 16304 15929 16313 15963
rect 16313 15929 16347 15963
rect 16347 15929 16356 15963
rect 16304 15920 16356 15929
rect 20352 15920 20404 15972
rect 20444 15920 20496 15972
rect 21088 15920 21140 15972
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 21456 15852 21508 15904
rect 24400 15895 24452 15904
rect 24400 15861 24409 15895
rect 24409 15861 24443 15895
rect 24443 15861 24452 15895
rect 24400 15852 24452 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 5724 15648 5776 15700
rect 5632 15512 5684 15564
rect 6736 15512 6788 15564
rect 7656 15648 7708 15700
rect 11520 15648 11572 15700
rect 12072 15648 12124 15700
rect 22284 15648 22336 15700
rect 15016 15580 15068 15632
rect 18512 15580 18564 15632
rect 20996 15580 21048 15632
rect 23940 15580 23992 15632
rect 18420 15512 18472 15564
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 20444 15512 20496 15564
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17776 15444 17828 15496
rect 21824 15512 21876 15564
rect 22100 15512 22152 15564
rect 24860 15512 24912 15564
rect 6920 15376 6972 15428
rect 11060 15376 11112 15428
rect 17408 15376 17460 15428
rect 20168 15376 20220 15428
rect 20812 15376 20864 15428
rect 24400 15376 24452 15428
rect 9404 15308 9456 15360
rect 14464 15351 14516 15360
rect 14464 15317 14473 15351
rect 14473 15317 14507 15351
rect 14507 15317 14516 15351
rect 14464 15308 14516 15317
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 18880 15308 18932 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 7564 15147 7616 15156
rect 7564 15113 7573 15147
rect 7573 15113 7607 15147
rect 7607 15113 7616 15147
rect 7564 15104 7616 15113
rect 9128 15104 9180 15156
rect 7840 15036 7892 15088
rect 9680 15104 9732 15156
rect 10048 15104 10100 15156
rect 11060 15104 11112 15156
rect 12808 15104 12860 15156
rect 14832 15104 14884 15156
rect 19064 15104 19116 15156
rect 19524 15104 19576 15156
rect 6920 14968 6972 15020
rect 12440 15079 12492 15088
rect 12440 15045 12449 15079
rect 12449 15045 12483 15079
rect 12483 15045 12492 15079
rect 12440 15036 12492 15045
rect 13636 15036 13688 15088
rect 15292 15036 15344 15088
rect 15844 15036 15896 15088
rect 24860 15036 24912 15088
rect 8576 14900 8628 14952
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 9772 14900 9824 14952
rect 12440 14832 12492 14884
rect 13360 14968 13412 15020
rect 13452 14968 13504 15020
rect 18512 14968 18564 15020
rect 21180 14968 21232 15020
rect 22192 15011 22244 15020
rect 22192 14977 22201 15011
rect 22201 14977 22235 15011
rect 22235 14977 22244 15011
rect 22192 14968 22244 14977
rect 24216 14968 24268 15020
rect 12808 14900 12860 14952
rect 13544 14900 13596 14952
rect 14096 14900 14148 14952
rect 13268 14832 13320 14884
rect 17224 14832 17276 14884
rect 22468 14900 22520 14952
rect 24768 14943 24820 14952
rect 24768 14909 24777 14943
rect 24777 14909 24811 14943
rect 24811 14909 24820 14943
rect 24768 14900 24820 14909
rect 10324 14764 10376 14816
rect 11428 14764 11480 14816
rect 13360 14764 13412 14816
rect 13544 14764 13596 14816
rect 18328 14764 18380 14816
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 9588 14560 9640 14612
rect 10508 14560 10560 14612
rect 11796 14560 11848 14612
rect 17132 14560 17184 14612
rect 12624 14492 12676 14544
rect 8760 14424 8812 14476
rect 9036 14424 9088 14476
rect 12808 14424 12860 14476
rect 14280 14424 14332 14476
rect 16856 14424 16908 14476
rect 9404 14356 9456 14408
rect 10232 14356 10284 14408
rect 13084 14356 13136 14408
rect 13912 14356 13964 14408
rect 14832 14356 14884 14408
rect 18604 14356 18656 14408
rect 20628 14399 20680 14408
rect 20628 14365 20637 14399
rect 20637 14365 20671 14399
rect 20671 14365 20680 14399
rect 20628 14356 20680 14365
rect 22376 14356 22428 14408
rect 7196 14288 7248 14340
rect 7564 14288 7616 14340
rect 10324 14288 10376 14340
rect 11152 14288 11204 14340
rect 13452 14288 13504 14340
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 16028 14288 16080 14340
rect 17960 14288 18012 14340
rect 21272 14288 21324 14340
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 9036 14220 9088 14272
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 12348 14220 12400 14272
rect 17408 14220 17460 14272
rect 20076 14220 20128 14272
rect 23388 14220 23440 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9220 14016 9272 14068
rect 9496 14016 9548 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13452 14016 13504 14068
rect 17316 14016 17368 14068
rect 8576 13948 8628 14000
rect 10140 13948 10192 14000
rect 10784 13948 10836 14000
rect 15568 13948 15620 14000
rect 15660 13948 15712 14000
rect 16028 13948 16080 14000
rect 18420 14016 18472 14068
rect 18696 14016 18748 14068
rect 20996 14016 21048 14068
rect 24584 14016 24636 14068
rect 19800 13948 19852 14000
rect 23296 13948 23348 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 2596 13880 2648 13932
rect 8760 13880 8812 13932
rect 10508 13880 10560 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 11980 13880 12032 13932
rect 13452 13880 13504 13932
rect 14096 13880 14148 13932
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 18420 13880 18472 13932
rect 18788 13880 18840 13932
rect 21548 13880 21600 13932
rect 22284 13880 22336 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 12716 13812 12768 13864
rect 14372 13744 14424 13796
rect 16672 13812 16724 13864
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 20260 13744 20312 13796
rect 21456 13812 21508 13864
rect 23480 13880 23532 13932
rect 14556 13676 14608 13728
rect 18788 13676 18840 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 21272 13676 21324 13728
rect 21456 13676 21508 13728
rect 22652 13719 22704 13728
rect 22652 13685 22661 13719
rect 22661 13685 22695 13719
rect 22695 13685 22704 13719
rect 22652 13676 22704 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 13268 13472 13320 13524
rect 13544 13472 13596 13524
rect 21272 13472 21324 13524
rect 23296 13515 23348 13524
rect 23296 13481 23305 13515
rect 23305 13481 23339 13515
rect 23339 13481 23348 13515
rect 23296 13472 23348 13481
rect 13452 13404 13504 13456
rect 16028 13404 16080 13456
rect 18880 13404 18932 13456
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7748 13336 7800 13388
rect 11152 13336 11204 13388
rect 18328 13336 18380 13388
rect 18696 13379 18748 13388
rect 18696 13345 18705 13379
rect 18705 13345 18739 13379
rect 18739 13345 18748 13379
rect 18696 13336 18748 13345
rect 20628 13336 20680 13388
rect 21640 13336 21692 13388
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 9036 13268 9088 13320
rect 13820 13268 13872 13320
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 17224 13268 17276 13320
rect 18788 13268 18840 13320
rect 19248 13268 19300 13320
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 7564 13200 7616 13252
rect 9680 13132 9732 13184
rect 16120 13200 16172 13252
rect 19616 13200 19668 13252
rect 20536 13200 20588 13252
rect 21088 13200 21140 13252
rect 21640 13200 21692 13252
rect 18512 13132 18564 13184
rect 20260 13132 20312 13184
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 9312 12928 9364 12980
rect 11704 12928 11756 12980
rect 15292 12928 15344 12980
rect 12808 12860 12860 12912
rect 13360 12860 13412 12912
rect 14556 12903 14608 12912
rect 14556 12869 14565 12903
rect 14565 12869 14599 12903
rect 14599 12869 14608 12903
rect 14556 12860 14608 12869
rect 6552 12792 6604 12844
rect 13544 12792 13596 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 15660 12792 15712 12844
rect 9680 12724 9732 12776
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 17316 12971 17368 12980
rect 17316 12937 17325 12971
rect 17325 12937 17359 12971
rect 17359 12937 17368 12971
rect 17316 12928 17368 12937
rect 18512 12971 18564 12980
rect 18512 12937 18521 12971
rect 18521 12937 18555 12971
rect 18555 12937 18564 12971
rect 18512 12928 18564 12937
rect 18328 12860 18380 12912
rect 16212 12792 16264 12844
rect 20260 12860 20312 12912
rect 20628 12860 20680 12912
rect 24860 12860 24912 12912
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22836 12792 22888 12844
rect 19248 12724 19300 12776
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 14280 12656 14332 12708
rect 19524 12656 19576 12708
rect 10968 12588 11020 12640
rect 19708 12588 19760 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 11152 12427 11204 12436
rect 11152 12393 11161 12427
rect 11161 12393 11195 12427
rect 11195 12393 11204 12427
rect 11152 12384 11204 12393
rect 13636 12384 13688 12436
rect 14924 12384 14976 12436
rect 16488 12384 16540 12436
rect 16580 12384 16632 12436
rect 22100 12384 22152 12436
rect 2780 12316 2832 12368
rect 4896 12316 4948 12368
rect 13452 12316 13504 12368
rect 14740 12316 14792 12368
rect 9680 12291 9732 12300
rect 9680 12257 9689 12291
rect 9689 12257 9723 12291
rect 9723 12257 9732 12291
rect 9680 12248 9732 12257
rect 10968 12248 11020 12300
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 11888 12180 11940 12232
rect 13636 12180 13688 12232
rect 13820 12248 13872 12300
rect 16396 12316 16448 12368
rect 20076 12316 20128 12368
rect 19340 12248 19392 12300
rect 20628 12248 20680 12300
rect 22376 12180 22428 12232
rect 24584 12180 24636 12232
rect 10140 12112 10192 12164
rect 13360 12112 13412 12164
rect 14740 12155 14792 12164
rect 14740 12121 14749 12155
rect 14749 12121 14783 12155
rect 14783 12121 14792 12155
rect 14740 12112 14792 12121
rect 15200 12112 15252 12164
rect 16764 12112 16816 12164
rect 12440 12044 12492 12096
rect 14372 12044 14424 12096
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 18696 12112 18748 12164
rect 19432 12112 19484 12164
rect 25320 12112 25372 12164
rect 18420 12044 18472 12096
rect 19616 12087 19668 12096
rect 19616 12053 19625 12087
rect 19625 12053 19659 12087
rect 19659 12053 19668 12087
rect 19616 12044 19668 12053
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 13820 11840 13872 11892
rect 14556 11840 14608 11892
rect 14924 11883 14976 11892
rect 14924 11849 14933 11883
rect 14933 11849 14967 11883
rect 14967 11849 14976 11883
rect 14924 11840 14976 11849
rect 15660 11772 15712 11824
rect 17132 11840 17184 11892
rect 9404 11636 9456 11688
rect 11244 11636 11296 11688
rect 14648 11704 14700 11756
rect 11980 11568 12032 11620
rect 15292 11636 15344 11688
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 16212 11568 16264 11620
rect 17408 11772 17460 11824
rect 19340 11772 19392 11824
rect 22376 11883 22428 11892
rect 22376 11849 22385 11883
rect 22385 11849 22419 11883
rect 22419 11849 22428 11883
rect 22376 11840 22428 11849
rect 16856 11704 16908 11756
rect 19524 11704 19576 11756
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 23848 11704 23900 11756
rect 19984 11636 20036 11688
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 19340 11568 19392 11620
rect 19800 11568 19852 11620
rect 22836 11568 22888 11620
rect 19432 11500 19484 11552
rect 23940 11500 23992 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 13820 11296 13872 11348
rect 22560 11296 22612 11348
rect 23296 11296 23348 11348
rect 10876 11228 10928 11280
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 13544 11228 13596 11280
rect 14372 11228 14424 11280
rect 15752 11092 15804 11144
rect 16396 11092 16448 11144
rect 22192 11228 22244 11280
rect 19708 11160 19760 11212
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 20720 11160 20772 11212
rect 22652 11160 22704 11212
rect 10140 11024 10192 11076
rect 11152 11024 11204 11076
rect 11980 11024 12032 11076
rect 12808 11024 12860 11076
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 15016 10956 15068 11008
rect 16028 11024 16080 11076
rect 23388 11024 23440 11076
rect 22744 10999 22796 11008
rect 22744 10965 22753 10999
rect 22753 10965 22787 10999
rect 22787 10965 22796 10999
rect 22744 10956 22796 10965
rect 23848 10999 23900 11008
rect 23848 10965 23857 10999
rect 23857 10965 23891 10999
rect 23891 10965 23900 10999
rect 23848 10956 23900 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 19248 10752 19300 10804
rect 19984 10752 20036 10804
rect 18328 10727 18380 10736
rect 18328 10693 18337 10727
rect 18337 10693 18371 10727
rect 18371 10693 18380 10727
rect 18328 10684 18380 10693
rect 19432 10616 19484 10668
rect 19800 10616 19852 10668
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 24676 10412 24728 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 23756 10072 23808 10124
rect 9864 10004 9916 10056
rect 20168 10004 20220 10056
rect 24584 10004 24636 10056
rect 24952 9936 25004 9988
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 14832 9868 14884 9920
rect 24584 9911 24636 9920
rect 24584 9877 24593 9911
rect 24593 9877 24627 9911
rect 24627 9877 24636 9911
rect 24584 9868 24636 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 14188 9596 14240 9648
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 23572 9528 23624 9580
rect 5540 9460 5592 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 15200 9392 15252 9444
rect 24032 9324 24084 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 3056 9120 3108 9172
rect 5908 9120 5960 9172
rect 22744 8984 22796 9036
rect 15936 8916 15988 8968
rect 18788 8916 18840 8968
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 17776 8848 17828 8900
rect 20720 8848 20772 8900
rect 5816 8780 5868 8832
rect 7564 8780 7616 8832
rect 22836 8780 22888 8832
rect 24124 8780 24176 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 6828 8576 6880 8628
rect 15752 8576 15804 8628
rect 16028 8576 16080 8628
rect 5816 8508 5868 8560
rect 12716 8508 12768 8560
rect 24860 8508 24912 8560
rect 25136 8551 25188 8560
rect 25136 8517 25145 8551
rect 25145 8517 25179 8551
rect 25179 8517 25188 8551
rect 25136 8508 25188 8517
rect 23848 8440 23900 8492
rect 2780 8372 2832 8424
rect 24492 8372 24544 8424
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 16580 7828 16632 7880
rect 20812 7828 20864 7880
rect 23296 7828 23348 7880
rect 24676 7828 24728 7880
rect 21272 7760 21324 7812
rect 24952 7760 25004 7812
rect 20444 7692 20496 7744
rect 24676 7735 24728 7744
rect 24676 7701 24685 7735
rect 24685 7701 24719 7735
rect 24719 7701 24728 7735
rect 24676 7692 24728 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 25412 7420 25464 7472
rect 20812 7352 20864 7404
rect 20904 7352 20956 7404
rect 24584 7352 24636 7404
rect 22468 7284 22520 7336
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 14556 6808 14608 6860
rect 16028 6740 16080 6792
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 19708 6672 19760 6724
rect 3148 6604 3200 6656
rect 6276 6604 6328 6656
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 24952 6740 25004 6792
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 23480 6672 23532 6724
rect 24492 6672 24544 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 20904 6400 20956 6452
rect 12072 6332 12124 6384
rect 17316 6264 17368 6316
rect 22376 6332 22428 6384
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 5172 6196 5224 6248
rect 11244 6196 11296 6248
rect 22192 6196 22244 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 20812 6060 20864 6112
rect 24768 6060 24820 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 22100 5856 22152 5908
rect 24768 5899 24820 5908
rect 24768 5865 24777 5899
rect 24777 5865 24811 5899
rect 24811 5865 24820 5899
rect 24768 5856 24820 5865
rect 20444 5788 20496 5840
rect 20628 5720 20680 5772
rect 2044 5652 2096 5704
rect 8484 5652 8536 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 10600 5584 10652 5636
rect 15844 5584 15896 5636
rect 21732 5584 21784 5636
rect 24492 5584 24544 5636
rect 2136 5516 2188 5568
rect 6460 5516 6512 5568
rect 9588 5516 9640 5568
rect 10324 5516 10376 5568
rect 22744 5516 22796 5568
rect 23848 5516 23900 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 18052 5176 18104 5228
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 19708 5176 19760 5228
rect 24676 5176 24728 5228
rect 19432 5108 19484 5160
rect 19524 5108 19576 5160
rect 22284 5108 22336 5160
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 9404 4972 9456 5024
rect 12624 4972 12676 5024
rect 23572 4972 23624 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 3240 4768 3292 4820
rect 6368 4768 6420 4820
rect 6460 4768 6512 4820
rect 11612 4768 11664 4820
rect 25320 4811 25372 4820
rect 25320 4777 25329 4811
rect 25329 4777 25363 4811
rect 25363 4777 25372 4811
rect 25320 4768 25372 4777
rect 18052 4632 18104 4684
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 19340 4564 19392 4616
rect 20536 4564 20588 4616
rect 18328 4539 18380 4548
rect 18328 4505 18337 4539
rect 18337 4505 18371 4539
rect 18371 4505 18380 4539
rect 18328 4496 18380 4505
rect 20352 4539 20404 4548
rect 20352 4505 20361 4539
rect 20361 4505 20395 4539
rect 20395 4505 20404 4539
rect 20352 4496 20404 4505
rect 21088 4496 21140 4548
rect 19800 4428 19852 4480
rect 23756 4564 23808 4616
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 5080 4156 5132 4208
rect 8944 4156 8996 4208
rect 11520 4156 11572 4208
rect 13728 4156 13780 4208
rect 21548 4156 21600 4208
rect 1124 4088 1176 4140
rect 8852 4088 8904 4140
rect 9220 4088 9272 4140
rect 13636 4088 13688 4140
rect 15200 4088 15252 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 12808 4020 12860 4072
rect 16212 4020 16264 4072
rect 18420 4020 18472 4072
rect 20260 4020 20312 4072
rect 5540 3952 5592 4004
rect 7840 3952 7892 4004
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 21548 3952 21600 4004
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 2780 3680 2832 3732
rect 3424 3680 3476 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 6736 3680 6788 3732
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 9588 3680 9640 3732
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 4988 3612 5040 3664
rect 16028 3612 16080 3664
rect 12532 3544 12584 3596
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 21364 3544 21416 3596
rect 23296 3544 23348 3596
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 2780 3476 2832 3528
rect 2872 3476 2924 3528
rect 4804 3476 4856 3528
rect 5540 3476 5592 3528
rect 6276 3476 6328 3528
rect 7380 3476 7432 3528
rect 7840 3476 7892 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 1492 3408 1544 3460
rect 10692 3476 10744 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 17776 3476 17828 3528
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 14464 3408 14516 3460
rect 19156 3408 19208 3460
rect 24308 3408 24360 3460
rect 14740 3340 14792 3392
rect 22008 3340 22060 3392
rect 22836 3340 22888 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 23756 3136 23808 3188
rect 3884 3068 3936 3120
rect 6092 3068 6144 3120
rect 1860 3000 1912 3052
rect 3332 3000 3384 3052
rect 3700 3000 3752 3052
rect 4436 3000 4488 3052
rect 5172 3000 5224 3052
rect 5908 3000 5960 3052
rect 15016 3068 15068 3120
rect 19432 3068 19484 3120
rect 23940 3068 23992 3120
rect 9404 3000 9456 3052
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12440 3000 12492 3052
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 16672 3000 16724 3052
rect 17868 3000 17920 3052
rect 23572 3043 23624 3052
rect 23572 3009 23581 3043
rect 23581 3009 23615 3043
rect 23615 3009 23624 3043
rect 23572 3000 23624 3009
rect 7012 2932 7064 2984
rect 8484 2932 8536 2984
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 11796 2932 11848 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 7288 2864 7340 2916
rect 16580 2864 16632 2916
rect 19892 2864 19944 2916
rect 21088 2864 21140 2916
rect 24492 2932 24544 2984
rect 25044 2864 25096 2916
rect 5080 2796 5132 2848
rect 9496 2796 9548 2848
rect 11060 2796 11112 2848
rect 17316 2796 17368 2848
rect 18328 2796 18380 2848
rect 18788 2796 18840 2848
rect 20352 2796 20404 2848
rect 20996 2796 21048 2848
rect 22284 2796 22336 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 2044 2635 2096 2644
rect 2044 2601 2053 2635
rect 2053 2601 2087 2635
rect 2087 2601 2096 2635
rect 2044 2592 2096 2601
rect 6460 2592 6512 2644
rect 10784 2592 10836 2644
rect 15292 2592 15344 2644
rect 8668 2524 8720 2576
rect 9496 2456 9548 2508
rect 2228 2388 2280 2440
rect 2596 2388 2648 2440
rect 4068 2388 4120 2440
rect 6644 2388 6696 2440
rect 15936 2524 15988 2576
rect 11704 2456 11756 2508
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 11428 2388 11480 2440
rect 14372 2456 14424 2508
rect 15108 2456 15160 2508
rect 16304 2388 16356 2440
rect 16764 2388 16816 2440
rect 16948 2388 17000 2440
rect 9036 2320 9088 2372
rect 12164 2320 12216 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 17040 2320 17092 2372
rect 21456 2388 21508 2440
rect 18512 2320 18564 2372
rect 7748 2252 7800 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 938 56200 994 57000
rect 1306 56200 1362 57000
rect 1674 56200 1730 57000
rect 2042 56200 2098 57000
rect 2410 56200 2466 57000
rect 2516 56222 2728 56250
rect 952 52630 980 56200
rect 1320 55214 1348 56200
rect 1228 55186 1348 55214
rect 940 52624 992 52630
rect 940 52566 992 52572
rect 940 50856 992 50862
rect 940 50798 992 50804
rect 952 50425 980 50798
rect 938 50416 994 50425
rect 938 50351 994 50360
rect 1228 49298 1256 55186
rect 1306 52728 1362 52737
rect 1306 52663 1362 52672
rect 1320 52562 1348 52663
rect 1308 52556 1360 52562
rect 1308 52498 1360 52504
rect 1688 49774 1716 56200
rect 2056 52698 2084 56200
rect 2424 56114 2452 56200
rect 2516 56114 2544 56222
rect 2424 56086 2544 56114
rect 2700 53122 2728 56222
rect 2778 56200 2834 57000
rect 3146 56200 3202 57000
rect 3514 56200 3570 57000
rect 3882 56200 3938 57000
rect 4250 56200 4306 57000
rect 4618 56200 4674 57000
rect 4986 56200 5042 57000
rect 5354 56200 5410 57000
rect 5722 56200 5778 57000
rect 6090 56200 6146 57000
rect 6458 56200 6514 57000
rect 6826 56200 6882 57000
rect 6932 56222 7144 56250
rect 2792 55214 2820 56200
rect 3160 55214 3188 56200
rect 2792 55186 2912 55214
rect 3160 55186 3372 55214
rect 2778 55040 2834 55049
rect 2778 54975 2834 54984
rect 2792 53242 2820 54975
rect 2780 53236 2832 53242
rect 2780 53178 2832 53184
rect 2700 53094 2820 53122
rect 2044 52692 2096 52698
rect 2044 52634 2096 52640
rect 2792 51474 2820 53094
rect 2780 51468 2832 51474
rect 2780 51410 2832 51416
rect 2884 50862 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 52494 3372 55186
rect 3424 52692 3476 52698
rect 3424 52634 3476 52640
rect 3148 52488 3200 52494
rect 3148 52430 3200 52436
rect 3332 52488 3384 52494
rect 3332 52430 3384 52436
rect 3160 52306 3188 52430
rect 3160 52278 3372 52306
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 50856 2924 50862
rect 2872 50798 2924 50804
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 1768 49836 1820 49842
rect 1768 49778 1820 49784
rect 1676 49768 1728 49774
rect 1676 49710 1728 49716
rect 1216 49292 1268 49298
rect 1216 49234 1268 49240
rect 1584 49224 1636 49230
rect 1584 49166 1636 49172
rect 938 48104 994 48113
rect 938 48039 940 48048
rect 992 48039 994 48048
rect 940 48010 992 48016
rect 940 45960 992 45966
rect 940 45902 992 45908
rect 952 45801 980 45902
rect 938 45792 994 45801
rect 938 45727 994 45736
rect 1596 40730 1624 49166
rect 1780 42362 1808 49778
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 3344 45554 3372 52278
rect 3436 50386 3464 52634
rect 3528 51950 3556 56200
rect 3896 53258 3924 56200
rect 3896 53230 4200 53258
rect 3976 52896 4028 52902
rect 3976 52838 4028 52844
rect 3516 51944 3568 51950
rect 3516 51886 3568 51892
rect 3700 50924 3752 50930
rect 3700 50866 3752 50872
rect 3424 50380 3476 50386
rect 3424 50322 3476 50328
rect 3516 50312 3568 50318
rect 3516 50254 3568 50260
rect 3344 45526 3464 45554
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 1768 42356 1820 42362
rect 1768 42298 1820 42304
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 3436 41818 3464 45526
rect 3424 41812 3476 41818
rect 3424 41754 3476 41760
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41177 1716 41482
rect 3528 41274 3556 50254
rect 3712 42770 3740 50866
rect 3988 48822 4016 52838
rect 4172 51474 4200 53230
rect 4264 53174 4292 56200
rect 4632 53650 4660 56200
rect 4712 54188 4764 54194
rect 4712 54130 4764 54136
rect 4620 53644 4672 53650
rect 4620 53586 4672 53592
rect 4252 53168 4304 53174
rect 4252 53110 4304 53116
rect 4252 52896 4304 52902
rect 4252 52838 4304 52844
rect 4160 51468 4212 51474
rect 4160 51410 4212 51416
rect 4264 51406 4292 52838
rect 4436 52624 4488 52630
rect 4436 52566 4488 52572
rect 4252 51400 4304 51406
rect 4252 51342 4304 51348
rect 4448 50386 4476 52566
rect 4724 51610 4752 54130
rect 5000 51950 5028 56200
rect 5368 54262 5396 56200
rect 5356 54256 5408 54262
rect 5356 54198 5408 54204
rect 5448 53576 5500 53582
rect 5448 53518 5500 53524
rect 4988 51944 5040 51950
rect 4988 51886 5040 51892
rect 4712 51604 4764 51610
rect 4712 51546 4764 51552
rect 4436 50380 4488 50386
rect 4436 50322 4488 50328
rect 3976 48816 4028 48822
rect 3976 48758 4028 48764
rect 3884 48068 3936 48074
rect 3884 48010 3936 48016
rect 3700 42764 3752 42770
rect 3700 42706 3752 42712
rect 3792 42220 3844 42226
rect 3792 42162 3844 42168
rect 3516 41268 3568 41274
rect 3516 41210 3568 41216
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 1584 40724 1636 40730
rect 1584 40666 1636 40672
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 940 38956 992 38962
rect 940 38898 992 38904
rect 952 38865 980 38898
rect 938 38856 994 38865
rect 938 38791 994 38800
rect 1860 38752 1912 38758
rect 1860 38694 1912 38700
rect 940 36780 992 36786
rect 940 36722 992 36728
rect 952 36553 980 36722
rect 938 36544 994 36553
rect 938 36479 994 36488
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1780 34241 1808 34546
rect 1766 34232 1822 34241
rect 1766 34167 1822 34176
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 952 31929 980 32370
rect 1584 32224 1636 32230
rect 1584 32166 1636 32172
rect 938 31920 994 31929
rect 938 31855 994 31864
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1320 29617 1348 29650
rect 1306 29608 1362 29617
rect 1306 29543 1362 29552
rect 1308 27532 1360 27538
rect 1308 27474 1360 27480
rect 1320 27305 1348 27474
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1596 26450 1624 32166
rect 1872 29646 1900 38694
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 3424 36576 3476 36582
rect 3424 36518 3476 36524
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 3332 34740 3384 34746
rect 3332 34682 3384 34688
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1860 29640 1912 29646
rect 1860 29582 1912 29588
rect 1780 27130 1808 29582
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3344 27538 3372 34682
rect 3436 28626 3464 36518
rect 3804 31754 3832 42162
rect 3896 40050 3924 48010
rect 5460 45554 5488 53518
rect 5736 53174 5764 56200
rect 5724 53168 5776 53174
rect 5724 53110 5776 53116
rect 6104 52562 6132 56200
rect 6368 53100 6420 53106
rect 6368 53042 6420 53048
rect 6000 52556 6052 52562
rect 6000 52498 6052 52504
rect 6092 52556 6144 52562
rect 6092 52498 6144 52504
rect 5724 52488 5776 52494
rect 5724 52430 5776 52436
rect 5632 52080 5684 52086
rect 5632 52022 5684 52028
rect 5540 51264 5592 51270
rect 5540 51206 5592 51212
rect 5552 51066 5580 51206
rect 5540 51060 5592 51066
rect 5540 51002 5592 51008
rect 5540 50312 5592 50318
rect 5540 50254 5592 50260
rect 5368 45526 5488 45554
rect 5172 43308 5224 43314
rect 5172 43250 5224 43256
rect 4160 42628 4212 42634
rect 4160 42570 4212 42576
rect 3976 41540 4028 41546
rect 3976 41482 4028 41488
rect 3884 40044 3936 40050
rect 3884 39986 3936 39992
rect 3988 31754 4016 41482
rect 4172 41414 4200 42570
rect 4172 41386 4292 41414
rect 4068 41132 4120 41138
rect 4068 41074 4120 41080
rect 3620 31726 3832 31754
rect 3896 31726 4016 31754
rect 3620 30054 3648 31726
rect 3896 31090 3924 31726
rect 3712 31062 3924 31090
rect 3608 30048 3660 30054
rect 3608 29990 3660 29996
rect 3516 29572 3568 29578
rect 3516 29514 3568 29520
rect 3424 28620 3476 28626
rect 3424 28562 3476 28568
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 1952 27464 2004 27470
rect 1952 27406 2004 27412
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1584 26444 1636 26450
rect 1584 26386 1636 26392
rect 1308 25356 1360 25362
rect 1308 25298 1360 25304
rect 1320 24993 1348 25298
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1306 24984 1362 24993
rect 1306 24919 1362 24928
rect 1308 23180 1360 23186
rect 1308 23122 1360 23128
rect 1320 22681 1348 23122
rect 1780 22778 1808 25230
rect 1964 24682 1992 27406
rect 3528 27130 3556 29514
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 2884 25770 2912 26930
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 2872 25764 2924 25770
rect 2872 25706 2924 25712
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 1952 24676 2004 24682
rect 1952 24618 2004 24624
rect 2228 24132 2280 24138
rect 2228 24074 2280 24080
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1306 22672 1362 22681
rect 1306 22607 1362 22616
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 20466 1808 21830
rect 2240 21486 2268 24074
rect 2792 23882 2820 24686
rect 2700 23866 2820 23882
rect 2688 23860 2820 23866
rect 2740 23854 2820 23860
rect 2688 23802 2740 23808
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2700 22234 2728 23054
rect 2884 22778 2912 24754
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 3344 23322 3372 25842
rect 3436 24070 3464 25842
rect 3620 25838 3648 26930
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3620 25158 3648 25774
rect 3712 25294 3740 31062
rect 4080 28422 4108 41074
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4172 34746 4200 35430
rect 4160 34740 4212 34746
rect 4160 34682 4212 34688
rect 4160 34400 4212 34406
rect 4160 34342 4212 34348
rect 4172 34202 4200 34342
rect 4160 34196 4212 34202
rect 4160 34138 4212 34144
rect 4264 31754 4292 41386
rect 5080 40452 5132 40458
rect 5080 40394 5132 40400
rect 4528 37800 4580 37806
rect 4528 37742 4580 37748
rect 4540 36650 4568 37742
rect 4988 37664 5040 37670
rect 4988 37606 5040 37612
rect 5000 37262 5028 37606
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4528 36644 4580 36650
rect 4528 36586 4580 36592
rect 4172 31726 4292 31754
rect 4172 31346 4200 31726
rect 4632 31482 4660 36722
rect 5000 36174 5028 37198
rect 4988 36168 5040 36174
rect 4988 36110 5040 36116
rect 5000 35494 5028 36110
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 5000 35086 5028 35430
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 4896 33992 4948 33998
rect 5000 33980 5028 35022
rect 4948 33952 5028 33980
rect 4896 33934 4948 33940
rect 4908 32978 4936 33934
rect 4896 32972 4948 32978
rect 4896 32914 4948 32920
rect 4908 31890 4936 32914
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4712 31816 4764 31822
rect 4712 31758 4764 31764
rect 4724 31482 4752 31758
rect 4620 31476 4672 31482
rect 4620 31418 4672 31424
rect 4712 31476 4764 31482
rect 4712 31418 4764 31424
rect 5092 31414 5120 40394
rect 5184 36922 5212 43250
rect 5368 42702 5396 45526
rect 5552 43450 5580 50254
rect 5540 43444 5592 43450
rect 5540 43386 5592 43392
rect 5356 42696 5408 42702
rect 5356 42638 5408 42644
rect 5644 41750 5672 52022
rect 5736 46170 5764 52430
rect 5724 46164 5776 46170
rect 5724 46106 5776 46112
rect 6012 45554 6040 52498
rect 6276 52012 6328 52018
rect 6276 51954 6328 51960
rect 6012 45526 6132 45554
rect 5632 41744 5684 41750
rect 5632 41686 5684 41692
rect 5356 41540 5408 41546
rect 5356 41482 5408 41488
rect 5368 41414 5396 41482
rect 5368 41386 5488 41414
rect 5172 36916 5224 36922
rect 5172 36858 5224 36864
rect 5264 36644 5316 36650
rect 5264 36586 5316 36592
rect 5276 34746 5304 36586
rect 5264 34740 5316 34746
rect 5264 34682 5316 34688
rect 5356 34196 5408 34202
rect 5356 34138 5408 34144
rect 5080 31408 5132 31414
rect 5080 31350 5132 31356
rect 4160 31340 4212 31346
rect 4160 31282 4212 31288
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 3884 26308 3936 26314
rect 3884 26250 3936 26256
rect 3792 25764 3844 25770
rect 3792 25706 3844 25712
rect 3700 25288 3752 25294
rect 3700 25230 3752 25236
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2792 21622 2820 22510
rect 2884 22114 2912 22578
rect 3436 22574 3464 24006
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2884 22086 3004 22114
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1308 20392 1360 20398
rect 1306 20360 1308 20369
rect 1360 20360 1362 20369
rect 1306 20295 1362 20304
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1320 18057 1348 18158
rect 1306 18048 1362 18057
rect 1306 17983 1362 17992
rect 1780 16114 1808 18566
rect 1872 18290 1900 19654
rect 2240 18766 2268 21422
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2792 21010 2820 21286
rect 2884 21146 2912 21966
rect 2976 21690 3004 22086
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 2884 16794 2912 20878
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19854 3372 21558
rect 3528 20942 3556 22578
rect 3620 22098 3648 25094
rect 3608 22092 3660 22098
rect 3804 22094 3832 25706
rect 3896 22778 3924 26250
rect 3988 26042 4016 28358
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3988 24614 4016 25230
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 4080 24410 4108 27270
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4908 26450 4936 26726
rect 4896 26444 4948 26450
rect 4896 26386 4948 26392
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4632 24614 4660 25434
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4080 23730 4108 23802
rect 4068 23724 4120 23730
rect 3988 23684 4068 23712
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3804 22066 3924 22094
rect 3608 22034 3660 22040
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3804 18970 3832 21490
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15745 1348 15982
rect 1306 15736 1362 15745
rect 1306 15671 1362 15680
rect 2608 13938 2636 16390
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13433 2820 13806
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2778 13424 2834 13433
rect 2778 13359 2834 13368
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2792 11121 2820 12310
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2778 11112 2834 11121
rect 2778 11047 2834 11056
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3068 8809 3096 9114
rect 3054 8800 3110 8809
rect 3054 8735 3110 8744
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1124 4140 1176 4146
rect 1124 4082 1176 4088
rect 1136 800 1164 4082
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1504 800 1532 3402
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 800 1900 2994
rect 2056 2650 2084 5646
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 3194 2176 5510
rect 2792 3738 2820 8366
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6497 3188 6598
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3252 4185 3280 4762
rect 3238 4176 3294 4185
rect 3238 4111 3294 4120
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3436 3738 3464 18770
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2240 800 2268 2382
rect 2608 800 2636 2382
rect 2792 1873 2820 3470
rect 2778 1864 2834 1873
rect 2884 1850 2912 3470
rect 3896 3126 3924 22066
rect 3988 21010 4016 23684
rect 4068 23666 4120 23672
rect 4264 23526 4292 24278
rect 4448 24274 4476 24550
rect 4436 24268 4488 24274
rect 4436 24210 4488 24216
rect 4252 23520 4304 23526
rect 4252 23462 4304 23468
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 4172 21554 4200 22374
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4264 21010 4292 23462
rect 4448 21554 4476 24210
rect 4632 23662 4660 24550
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 17338 4200 18702
rect 4448 17882 4476 21490
rect 4816 19514 4844 22442
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4908 12374 4936 26386
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 5000 23662 5028 23734
rect 4988 23656 5040 23662
rect 4988 23598 5040 23604
rect 5092 22094 5120 31350
rect 5368 31278 5396 34138
rect 5356 31272 5408 31278
rect 5356 31214 5408 31220
rect 5460 31210 5488 41386
rect 6104 40118 6132 45526
rect 6288 44538 6316 51954
rect 6380 45082 6408 53042
rect 6472 52494 6500 56200
rect 6840 55214 6868 56200
rect 6748 55186 6868 55214
rect 6644 53508 6696 53514
rect 6644 53450 6696 53456
rect 6552 53032 6604 53038
rect 6552 52974 6604 52980
rect 6460 52488 6512 52494
rect 6460 52430 6512 52436
rect 6564 52306 6592 52974
rect 6472 52278 6592 52306
rect 6368 45076 6420 45082
rect 6368 45018 6420 45024
rect 6276 44532 6328 44538
rect 6276 44474 6328 44480
rect 6472 42770 6500 52278
rect 6656 45554 6684 53450
rect 6748 53394 6776 55186
rect 6932 54346 6960 56222
rect 7116 56114 7144 56222
rect 7194 56200 7250 57000
rect 7562 56200 7618 57000
rect 7930 56200 7986 57000
rect 8298 56200 8354 57000
rect 8666 56200 8722 57000
rect 9034 56200 9090 57000
rect 9402 56200 9458 57000
rect 9770 56200 9826 57000
rect 10138 56200 10194 57000
rect 10506 56200 10562 57000
rect 10874 56200 10930 57000
rect 11242 56200 11298 57000
rect 11610 56200 11666 57000
rect 11978 56200 12034 57000
rect 12346 56200 12402 57000
rect 12714 56200 12770 57000
rect 13082 56200 13138 57000
rect 13188 56222 13400 56250
rect 7208 56114 7236 56200
rect 7116 56086 7236 56114
rect 6840 54318 6960 54346
rect 6840 54262 6868 54318
rect 6828 54256 6880 54262
rect 6828 54198 6880 54204
rect 7472 54188 7524 54194
rect 7472 54130 7524 54136
rect 7380 53576 7432 53582
rect 7380 53518 7432 53524
rect 6748 53366 7052 53394
rect 6828 53100 6880 53106
rect 6828 53042 6880 53048
rect 6840 47258 6868 53042
rect 6920 52488 6972 52494
rect 6920 52430 6972 52436
rect 6932 51474 6960 52430
rect 7024 51950 7052 53366
rect 7104 52012 7156 52018
rect 7104 51954 7156 51960
rect 7012 51944 7064 51950
rect 7012 51886 7064 51892
rect 6920 51468 6972 51474
rect 6920 51410 6972 51416
rect 7012 51332 7064 51338
rect 7012 51274 7064 51280
rect 6920 50312 6972 50318
rect 6920 50254 6972 50260
rect 6828 47252 6880 47258
rect 6828 47194 6880 47200
rect 6564 45526 6684 45554
rect 6564 43994 6592 45526
rect 6932 44266 6960 50254
rect 7024 46714 7052 51274
rect 7116 50522 7144 51954
rect 7288 51400 7340 51406
rect 7288 51342 7340 51348
rect 7196 50924 7248 50930
rect 7196 50866 7248 50872
rect 7104 50516 7156 50522
rect 7104 50458 7156 50464
rect 7104 49836 7156 49842
rect 7104 49778 7156 49784
rect 7012 46708 7064 46714
rect 7012 46650 7064 46656
rect 7116 45554 7144 49778
rect 7208 45558 7236 50866
rect 7300 49858 7328 51342
rect 7392 49978 7420 53518
rect 7380 49972 7432 49978
rect 7380 49914 7432 49920
rect 7300 49830 7420 49858
rect 7288 45892 7340 45898
rect 7288 45834 7340 45840
rect 7024 45526 7144 45554
rect 7196 45552 7248 45558
rect 6920 44260 6972 44266
rect 6920 44202 6972 44208
rect 6552 43988 6604 43994
rect 6552 43930 6604 43936
rect 6460 42764 6512 42770
rect 6460 42706 6512 42712
rect 6460 42628 6512 42634
rect 6460 42570 6512 42576
rect 6920 42628 6972 42634
rect 6920 42570 6972 42576
rect 6276 41608 6328 41614
rect 6276 41550 6328 41556
rect 6288 41414 6316 41550
rect 6472 41414 6500 42570
rect 6288 41386 6408 41414
rect 6472 41386 6776 41414
rect 6276 41064 6328 41070
rect 6276 41006 6328 41012
rect 6288 40526 6316 41006
rect 6276 40520 6328 40526
rect 6276 40462 6328 40468
rect 6092 40112 6144 40118
rect 6092 40054 6144 40060
rect 6288 38418 6316 40462
rect 6276 38412 6328 38418
rect 6276 38354 6328 38360
rect 5540 38276 5592 38282
rect 5540 38218 5592 38224
rect 5552 37942 5580 38218
rect 5540 37936 5592 37942
rect 5540 37878 5592 37884
rect 5552 37194 5580 37878
rect 6184 37460 6236 37466
rect 6184 37402 6236 37408
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5552 36038 5580 37130
rect 6092 36712 6144 36718
rect 6092 36654 6144 36660
rect 6104 36174 6132 36654
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5552 35766 5580 35974
rect 5540 35760 5592 35766
rect 5540 35702 5592 35708
rect 5552 35018 5580 35702
rect 5540 35012 5592 35018
rect 5540 34954 5592 34960
rect 5552 34678 5580 34954
rect 5540 34672 5592 34678
rect 5592 34620 5672 34626
rect 5540 34614 5672 34620
rect 5552 34598 5672 34614
rect 5644 33930 5672 34598
rect 5632 33924 5684 33930
rect 5632 33866 5684 33872
rect 5448 31204 5500 31210
rect 5448 31146 5500 31152
rect 6000 29572 6052 29578
rect 6000 29514 6052 29520
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5828 25498 5856 28426
rect 5908 27056 5960 27062
rect 5908 26998 5960 27004
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5552 23186 5580 23802
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5828 23322 5856 23462
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5724 23044 5776 23050
rect 5724 22986 5776 22992
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5644 22234 5672 22578
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5092 22066 5212 22094
rect 5184 17270 5212 22066
rect 5736 21690 5764 22986
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 5644 19786 5672 20810
rect 5736 20806 5764 21286
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5460 18766 5488 19654
rect 5644 19174 5672 19722
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5460 17746 5488 18702
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5184 12434 5212 17206
rect 5460 16946 5488 17682
rect 5460 16918 5672 16946
rect 5644 16590 5672 16918
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5644 15570 5672 16526
rect 5736 15706 5764 20742
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5092 12406 5212 12434
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5092 6914 5120 12406
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5000 6886 5120 6914
rect 5000 3670 5028 6886
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5092 3738 5120 4150
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2884 1822 3004 1850
rect 2778 1799 2834 1808
rect 2976 800 3004 1822
rect 3344 800 3372 2994
rect 3712 800 3740 2994
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 800 4108 2382
rect 4448 800 4476 2994
rect 4816 800 4844 3470
rect 5184 3194 5212 6190
rect 5552 4010 5580 9454
rect 5920 9178 5948 26998
rect 6012 24886 6040 29514
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 6104 27062 6132 27338
rect 6092 27056 6144 27062
rect 6092 26998 6144 27004
rect 6196 26234 6224 37402
rect 6380 31754 6408 41386
rect 6552 40452 6604 40458
rect 6552 40394 6604 40400
rect 6564 39846 6592 40394
rect 6552 39840 6604 39846
rect 6552 39782 6604 39788
rect 6564 38010 6592 39782
rect 6552 38004 6604 38010
rect 6552 37946 6604 37952
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 6564 32842 6592 34682
rect 6748 34202 6776 41386
rect 6932 39642 6960 42570
rect 7024 42566 7052 45526
rect 7196 45494 7248 45500
rect 7196 44396 7248 44402
rect 7196 44338 7248 44344
rect 7208 44305 7236 44338
rect 7194 44296 7250 44305
rect 7194 44231 7250 44240
rect 7104 42696 7156 42702
rect 7104 42638 7156 42644
rect 7012 42560 7064 42566
rect 7012 42502 7064 42508
rect 7012 41268 7064 41274
rect 7012 41210 7064 41216
rect 6920 39636 6972 39642
rect 6920 39578 6972 39584
rect 6920 39500 6972 39506
rect 6920 39442 6972 39448
rect 6932 38554 6960 39442
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 6932 37330 6960 38490
rect 7024 38010 7052 41210
rect 7012 38004 7064 38010
rect 7012 37946 7064 37952
rect 7024 37466 7052 37946
rect 7012 37460 7064 37466
rect 7012 37402 7064 37408
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 7012 37324 7064 37330
rect 7012 37266 7064 37272
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 6840 36106 6868 36790
rect 6828 36100 6880 36106
rect 6828 36042 6880 36048
rect 7024 35834 7052 37266
rect 7012 35828 7064 35834
rect 7012 35770 7064 35776
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 6840 35018 6868 35566
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6828 35012 6880 35018
rect 6828 34954 6880 34960
rect 6736 34196 6788 34202
rect 6736 34138 6788 34144
rect 6828 34060 6880 34066
rect 6828 34002 6880 34008
rect 6840 33046 6868 34002
rect 6828 33040 6880 33046
rect 6828 32982 6880 32988
rect 6552 32836 6604 32842
rect 6552 32778 6604 32784
rect 6564 31822 6592 32778
rect 6828 32768 6880 32774
rect 6932 32722 6960 35090
rect 7024 34678 7052 35770
rect 7116 35290 7144 42638
rect 7300 41414 7328 45834
rect 7392 43994 7420 49830
rect 7484 45422 7512 54130
rect 7576 53650 7604 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7564 53644 7616 53650
rect 7564 53586 7616 53592
rect 7852 52562 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8312 53650 8340 56200
rect 8576 54120 8628 54126
rect 8576 54062 8628 54068
rect 8300 53644 8352 53650
rect 8300 53586 8352 53592
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7840 52556 7892 52562
rect 7840 52498 7892 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8392 50924 8444 50930
rect 8392 50866 8444 50872
rect 7564 50788 7616 50794
rect 7564 50730 7616 50736
rect 7472 45416 7524 45422
rect 7472 45358 7524 45364
rect 7576 44962 7604 50730
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7840 46572 7892 46578
rect 7840 46514 7892 46520
rect 7656 45484 7708 45490
rect 7656 45426 7708 45432
rect 7484 44934 7604 44962
rect 7380 43988 7432 43994
rect 7380 43930 7432 43936
rect 7300 41386 7420 41414
rect 7288 39908 7340 39914
rect 7288 39850 7340 39856
rect 7196 39636 7248 39642
rect 7196 39578 7248 39584
rect 7208 36582 7236 39578
rect 7300 37262 7328 39850
rect 7392 38350 7420 41386
rect 7484 39438 7512 44934
rect 7564 44804 7616 44810
rect 7564 44746 7616 44752
rect 7576 41274 7604 44746
rect 7564 41268 7616 41274
rect 7564 41210 7616 41216
rect 7564 41064 7616 41070
rect 7564 41006 7616 41012
rect 7576 40390 7604 41006
rect 7564 40384 7616 40390
rect 7564 40326 7616 40332
rect 7472 39432 7524 39438
rect 7472 39374 7524 39380
rect 7576 38554 7604 40326
rect 7668 39642 7696 45426
rect 7748 44396 7800 44402
rect 7748 44338 7800 44344
rect 7656 39636 7708 39642
rect 7656 39578 7708 39584
rect 7656 39296 7708 39302
rect 7656 39238 7708 39244
rect 7564 38548 7616 38554
rect 7564 38490 7616 38496
rect 7564 38412 7616 38418
rect 7564 38354 7616 38360
rect 7380 38344 7432 38350
rect 7380 38286 7432 38292
rect 7576 37874 7604 38354
rect 7564 37868 7616 37874
rect 7564 37810 7616 37816
rect 7288 37256 7340 37262
rect 7288 37198 7340 37204
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7104 35284 7156 35290
rect 7104 35226 7156 35232
rect 7300 35222 7328 37198
rect 7564 36712 7616 36718
rect 7564 36654 7616 36660
rect 7576 36242 7604 36654
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7288 35216 7340 35222
rect 7288 35158 7340 35164
rect 7564 35216 7616 35222
rect 7564 35158 7616 35164
rect 7012 34672 7064 34678
rect 7012 34614 7064 34620
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 6880 32716 6960 32722
rect 6828 32710 6960 32716
rect 6840 32694 6960 32710
rect 6932 32026 6960 32694
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6288 31726 6408 31754
rect 6288 30802 6316 31726
rect 7024 31482 7052 33594
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7392 30938 7420 31282
rect 7576 31278 7604 35158
rect 7668 34746 7696 39238
rect 7760 37126 7788 44338
rect 7852 41818 7880 46514
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 8404 45354 8432 50866
rect 8588 45554 8616 54062
rect 8680 53038 8708 56200
rect 9048 53650 9076 56200
rect 9416 54262 9444 56200
rect 9404 54256 9456 54262
rect 9404 54198 9456 54204
rect 9036 53644 9088 53650
rect 9036 53586 9088 53592
rect 9680 53644 9732 53650
rect 9680 53586 9732 53592
rect 9220 53100 9272 53106
rect 9220 53042 9272 53048
rect 9404 53100 9456 53106
rect 9404 53042 9456 53048
rect 8668 53032 8720 53038
rect 8668 52974 8720 52980
rect 8944 52488 8996 52494
rect 8944 52430 8996 52436
rect 8588 45526 8708 45554
rect 8392 45348 8444 45354
rect 8392 45290 8444 45296
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 8680 44538 8708 45526
rect 8668 44532 8720 44538
rect 8668 44474 8720 44480
rect 8956 43994 8984 52430
rect 9128 52012 9180 52018
rect 9128 51954 9180 51960
rect 9140 45082 9168 51954
rect 9128 45076 9180 45082
rect 9128 45018 9180 45024
rect 9036 44396 9088 44402
rect 9036 44338 9088 44344
rect 8944 43988 8996 43994
rect 8944 43930 8996 43936
rect 8300 43716 8352 43722
rect 8300 43658 8352 43664
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 8312 41614 8340 43658
rect 8576 42628 8628 42634
rect 8576 42570 8628 42576
rect 8392 42288 8444 42294
rect 8392 42230 8444 42236
rect 8300 41608 8352 41614
rect 8300 41550 8352 41556
rect 7840 41472 7892 41478
rect 8404 41426 8432 42230
rect 8484 42152 8536 42158
rect 8484 42094 8536 42100
rect 8496 41682 8524 42094
rect 8484 41676 8536 41682
rect 8484 41618 8536 41624
rect 7840 41414 7892 41420
rect 7852 38554 7880 41414
rect 8312 41398 8432 41426
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 8312 41138 8340 41398
rect 8496 41274 8524 41618
rect 8484 41268 8536 41274
rect 8484 41210 8536 41216
rect 8300 41132 8352 41138
rect 8300 41074 8352 41080
rect 8312 40458 8340 41074
rect 8300 40452 8352 40458
rect 8300 40394 8352 40400
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7840 38548 7892 38554
rect 7840 38490 7892 38496
rect 8024 38344 8076 38350
rect 8024 38286 8076 38292
rect 8036 38214 8064 38286
rect 7840 38208 7892 38214
rect 7840 38150 7892 38156
rect 8024 38208 8076 38214
rect 8024 38150 8076 38156
rect 8392 38208 8444 38214
rect 8392 38150 8444 38156
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7852 36378 7880 38150
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8300 37936 8352 37942
rect 8300 37878 8352 37884
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 8312 36854 8340 37878
rect 8404 37398 8432 38150
rect 8392 37392 8444 37398
rect 8392 37334 8444 37340
rect 8300 36848 8352 36854
rect 8300 36790 8352 36796
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7852 35034 7880 36314
rect 8312 36038 8340 36790
rect 8588 36310 8616 42570
rect 9048 41414 9076 44338
rect 9232 43926 9260 53042
rect 9416 50454 9444 53042
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9404 50448 9456 50454
rect 9404 50390 9456 50396
rect 9600 49910 9628 52430
rect 9692 51950 9720 53586
rect 9784 52562 9812 56200
rect 9864 54188 9916 54194
rect 9864 54130 9916 54136
rect 9772 52556 9824 52562
rect 9772 52498 9824 52504
rect 9680 51944 9732 51950
rect 9680 51886 9732 51892
rect 9876 51066 9904 54130
rect 10048 53576 10100 53582
rect 10048 53518 10100 53524
rect 9864 51060 9916 51066
rect 9864 51002 9916 51008
rect 9956 50924 10008 50930
rect 9956 50866 10008 50872
rect 9588 49904 9640 49910
rect 9588 49846 9640 49852
rect 9312 49836 9364 49842
rect 9312 49778 9364 49784
rect 9220 43920 9272 43926
rect 9220 43862 9272 43868
rect 9324 42566 9352 49778
rect 9772 48680 9824 48686
rect 9772 48622 9824 48628
rect 9404 48544 9456 48550
rect 9404 48486 9456 48492
rect 9416 44402 9444 48486
rect 9680 45960 9732 45966
rect 9680 45902 9732 45908
rect 9404 44396 9456 44402
rect 9404 44338 9456 44344
rect 9312 42560 9364 42566
rect 9312 42502 9364 42508
rect 9416 42022 9444 44338
rect 9496 43376 9548 43382
rect 9496 43318 9548 43324
rect 9508 43110 9536 43318
rect 9496 43104 9548 43110
rect 9496 43046 9548 43052
rect 9508 42362 9536 43046
rect 9496 42356 9548 42362
rect 9496 42298 9548 42304
rect 9404 42016 9456 42022
rect 9404 41958 9456 41964
rect 8864 41386 9076 41414
rect 8760 40180 8812 40186
rect 8760 40122 8812 40128
rect 8668 38752 8720 38758
rect 8668 38694 8720 38700
rect 8680 38350 8708 38694
rect 8668 38344 8720 38350
rect 8668 38286 8720 38292
rect 8772 37262 8800 40122
rect 8760 37256 8812 37262
rect 8760 37198 8812 37204
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 8760 36304 8812 36310
rect 8760 36246 8812 36252
rect 8300 36032 8352 36038
rect 8300 35974 8352 35980
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8312 35170 8340 35974
rect 8312 35142 8616 35170
rect 7852 35006 8340 35034
rect 7840 34944 7892 34950
rect 7840 34886 7892 34892
rect 7656 34740 7708 34746
rect 7656 34682 7708 34688
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7668 32314 7696 34478
rect 7748 34400 7800 34406
rect 7748 34342 7800 34348
rect 7760 33454 7788 34342
rect 7748 33448 7800 33454
rect 7748 33390 7800 33396
rect 7760 32978 7788 33390
rect 7748 32972 7800 32978
rect 7748 32914 7800 32920
rect 7760 32434 7788 32914
rect 7748 32428 7800 32434
rect 7748 32370 7800 32376
rect 7668 32286 7788 32314
rect 7656 32224 7708 32230
rect 7656 32166 7708 32172
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 7380 30932 7432 30938
rect 7380 30874 7432 30880
rect 6276 30796 6328 30802
rect 6276 30738 6328 30744
rect 7196 30796 7248 30802
rect 7196 30738 7248 30744
rect 6920 28620 6972 28626
rect 6920 28562 6972 28568
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6288 28014 6316 28494
rect 6276 28008 6328 28014
rect 6276 27950 6328 27956
rect 6288 27470 6316 27950
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 6288 26382 6316 27406
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6460 26308 6512 26314
rect 6460 26250 6512 26256
rect 6104 26206 6224 26234
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 23866 6040 24686
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6012 22574 6040 23802
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8566 5856 8774
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5078 2952 5134 2961
rect 5078 2887 5134 2896
rect 5092 2854 5120 2887
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5184 800 5212 2994
rect 5552 800 5580 3470
rect 6104 3126 6132 26206
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6184 24880 6236 24886
rect 6184 24822 6236 24828
rect 6196 21350 6224 24822
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 20806 6224 21286
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6196 19174 6224 19722
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18698 6224 19110
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6196 18358 6224 18634
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 6196 17678 6224 18294
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6196 16522 6224 17614
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 6288 6662 6316 25434
rect 6472 25362 6500 26250
rect 6932 25906 6960 28562
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6460 25356 6512 25362
rect 6460 25298 6512 25304
rect 6472 24750 6500 25298
rect 7024 24954 7052 26726
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7116 25362 7144 26522
rect 7208 25838 7236 30738
rect 7484 28914 7512 31214
rect 7576 29782 7604 31214
rect 7668 30734 7696 32166
rect 7760 30870 7788 32286
rect 7852 32026 7880 34886
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8312 34474 8340 35006
rect 8300 34468 8352 34474
rect 8300 34410 8352 34416
rect 8484 34400 8536 34406
rect 8484 34342 8536 34348
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 8404 31890 8432 32846
rect 8496 31890 8524 34342
rect 8588 33590 8616 35142
rect 8576 33584 8628 33590
rect 8576 33526 8628 33532
rect 8588 32570 8616 33526
rect 8668 32836 8720 32842
rect 8668 32778 8720 32784
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8680 32366 8708 32778
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 8404 31754 8432 31826
rect 8772 31754 8800 36246
rect 8312 31726 8432 31754
rect 8588 31726 8800 31754
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7852 31346 7880 31622
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 7748 30864 7800 30870
rect 7748 30806 7800 30812
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8312 30274 8340 31726
rect 8312 30246 8432 30274
rect 8404 30190 8432 30246
rect 8024 30184 8076 30190
rect 8024 30126 8076 30132
rect 8392 30184 8444 30190
rect 8392 30126 8444 30132
rect 7564 29776 7616 29782
rect 7564 29718 7616 29724
rect 8036 29714 8064 30126
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 7392 28886 7512 28914
rect 7288 28484 7340 28490
rect 7288 28426 7340 28432
rect 7300 28150 7328 28426
rect 7288 28144 7340 28150
rect 7288 28086 7340 28092
rect 7300 27402 7328 28086
rect 7288 27396 7340 27402
rect 7288 27338 7340 27344
rect 7300 26790 7328 27338
rect 7392 26926 7420 28886
rect 8220 28626 8248 29242
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 7300 26314 7328 26726
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 7196 25832 7248 25838
rect 7196 25774 7248 25780
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21146 6592 21830
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6380 4826 6408 20742
rect 6472 5574 6500 20742
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6564 17134 6592 17478
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16658 6592 17070
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 9450 6592 12786
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6656 6914 6684 23734
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6840 22166 6868 23258
rect 7024 23186 7052 24686
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 7116 23050 7144 23666
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7116 22216 7144 22986
rect 7024 22188 7144 22216
rect 6828 22160 6880 22166
rect 7024 22114 7052 22188
rect 6828 22102 6880 22108
rect 6932 22086 7052 22114
rect 7104 22092 7156 22098
rect 6932 22012 6960 22086
rect 7104 22034 7156 22040
rect 6840 21984 6960 22012
rect 7012 22024 7064 22030
rect 6840 20534 6868 21984
rect 7012 21966 7064 21972
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6840 19786 6868 20470
rect 7024 20058 7052 21966
rect 7116 20466 7144 22034
rect 7208 21570 7236 25638
rect 7392 22098 7420 26862
rect 7576 26586 7604 27814
rect 7852 27674 7880 28154
rect 8312 28014 8340 28358
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 7840 27668 7892 27674
rect 7840 27610 7892 27616
rect 7852 26858 7880 27610
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 8312 26926 8340 27950
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 7748 26852 7800 26858
rect 7748 26794 7800 26800
rect 7840 26852 7892 26858
rect 7840 26794 7892 26800
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7760 26518 7788 26794
rect 7748 26512 7800 26518
rect 7748 26454 7800 26460
rect 8404 26382 8432 27270
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 8404 25838 8432 26318
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7484 24274 7512 25298
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7852 24954 7880 25230
rect 8208 25152 8260 25158
rect 8260 25112 8340 25140
rect 8208 25094 8260 25100
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 8312 24834 8340 25112
rect 8220 24806 8340 24834
rect 8220 24750 8248 24806
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 8220 24206 8248 24550
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8496 24138 8524 29990
rect 8588 28626 8616 31726
rect 8864 29578 8892 41386
rect 9416 41070 9444 41958
rect 9588 41472 9640 41478
rect 9588 41414 9640 41420
rect 9404 41064 9456 41070
rect 9404 41006 9456 41012
rect 9416 40118 9444 41006
rect 9404 40112 9456 40118
rect 9404 40054 9456 40060
rect 9036 39500 9088 39506
rect 9036 39442 9088 39448
rect 9048 37738 9076 39442
rect 9496 39432 9548 39438
rect 9496 39374 9548 39380
rect 9404 39296 9456 39302
rect 9404 39238 9456 39244
rect 9312 38888 9364 38894
rect 9312 38830 9364 38836
rect 9324 37806 9352 38830
rect 9416 38554 9444 39238
rect 9508 38826 9536 39374
rect 9496 38820 9548 38826
rect 9496 38762 9548 38768
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 9600 38350 9628 41414
rect 9692 39370 9720 45902
rect 9784 44334 9812 48622
rect 9864 45960 9916 45966
rect 9864 45902 9916 45908
rect 9772 44328 9824 44334
rect 9772 44270 9824 44276
rect 9772 44192 9824 44198
rect 9772 44134 9824 44140
rect 9680 39364 9732 39370
rect 9680 39306 9732 39312
rect 9784 39098 9812 44134
rect 9876 42786 9904 45902
rect 9968 45354 9996 50866
rect 10060 45554 10088 53518
rect 10152 53038 10180 56200
rect 10520 53650 10548 56200
rect 10888 54262 10916 56200
rect 10876 54256 10928 54262
rect 10876 54198 10928 54204
rect 10508 53644 10560 53650
rect 10508 53586 10560 53592
rect 10508 53100 10560 53106
rect 10508 53042 10560 53048
rect 10140 53032 10192 53038
rect 10140 52974 10192 52980
rect 10520 51066 10548 53042
rect 11256 53038 11284 56200
rect 11624 53650 11652 56200
rect 11992 54126 12020 56200
rect 12072 54188 12124 54194
rect 12072 54130 12124 54136
rect 11980 54120 12032 54126
rect 11980 54062 12032 54068
rect 11612 53644 11664 53650
rect 11612 53586 11664 53592
rect 11704 53576 11756 53582
rect 11704 53518 11756 53524
rect 11244 53032 11296 53038
rect 11244 52974 11296 52980
rect 11716 52154 11744 53518
rect 12084 52698 12112 54130
rect 12072 52692 12124 52698
rect 12072 52634 12124 52640
rect 12360 52494 12388 56200
rect 12532 53440 12584 53446
rect 12532 53382 12584 53388
rect 11980 52488 12032 52494
rect 11980 52430 12032 52436
rect 12348 52488 12400 52494
rect 12348 52430 12400 52436
rect 11704 52148 11756 52154
rect 11704 52090 11756 52096
rect 11888 52012 11940 52018
rect 11888 51954 11940 51960
rect 10508 51060 10560 51066
rect 10508 51002 10560 51008
rect 10416 50244 10468 50250
rect 10416 50186 10468 50192
rect 10060 45526 10180 45554
rect 9956 45348 10008 45354
rect 9956 45290 10008 45296
rect 9956 44736 10008 44742
rect 9956 44678 10008 44684
rect 9968 44470 9996 44678
rect 9956 44464 10008 44470
rect 9956 44406 10008 44412
rect 9968 43654 9996 44406
rect 10152 44334 10180 45526
rect 10232 45484 10284 45490
rect 10232 45426 10284 45432
rect 10048 44328 10100 44334
rect 10048 44270 10100 44276
rect 10140 44328 10192 44334
rect 10140 44270 10192 44276
rect 10060 44180 10088 44270
rect 10244 44198 10272 45426
rect 10232 44192 10284 44198
rect 10060 44152 10180 44180
rect 9956 43648 10008 43654
rect 9956 43590 10008 43596
rect 9968 43110 9996 43590
rect 10048 43240 10100 43246
rect 10048 43182 10100 43188
rect 9956 43104 10008 43110
rect 9956 43046 10008 43052
rect 9876 42758 9996 42786
rect 9864 42696 9916 42702
rect 9864 42638 9916 42644
rect 9876 40050 9904 42638
rect 9968 42566 9996 42758
rect 10060 42634 10088 43182
rect 10152 42786 10180 44152
rect 10232 44134 10284 44140
rect 10324 43784 10376 43790
rect 10324 43726 10376 43732
rect 10232 43716 10284 43722
rect 10232 43658 10284 43664
rect 10244 42945 10272 43658
rect 10230 42936 10286 42945
rect 10230 42871 10286 42880
rect 10232 42832 10284 42838
rect 10152 42780 10232 42786
rect 10152 42774 10284 42780
rect 10152 42758 10272 42774
rect 10048 42628 10100 42634
rect 10048 42570 10100 42576
rect 9956 42560 10008 42566
rect 9956 42502 10008 42508
rect 10140 42560 10192 42566
rect 10140 42502 10192 42508
rect 9864 40044 9916 40050
rect 9864 39986 9916 39992
rect 9876 39914 9904 39986
rect 9864 39908 9916 39914
rect 9864 39850 9916 39856
rect 9864 39568 9916 39574
rect 9864 39510 9916 39516
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9876 38434 9904 39510
rect 10048 38956 10100 38962
rect 10048 38898 10100 38904
rect 9784 38406 9904 38434
rect 9588 38344 9640 38350
rect 9588 38286 9640 38292
rect 9784 38282 9812 38406
rect 9772 38276 9824 38282
rect 9772 38218 9824 38224
rect 9312 37800 9364 37806
rect 9312 37742 9364 37748
rect 9036 37732 9088 37738
rect 9036 37674 9088 37680
rect 9048 36378 9076 37674
rect 9324 36922 9352 37742
rect 9864 37188 9916 37194
rect 9864 37130 9916 37136
rect 9128 36916 9180 36922
rect 9128 36858 9180 36864
rect 9312 36916 9364 36922
rect 9312 36858 9364 36864
rect 9036 36372 9088 36378
rect 9036 36314 9088 36320
rect 9048 36145 9076 36314
rect 9034 36136 9090 36145
rect 9034 36071 9090 36080
rect 9048 31929 9076 36071
rect 9140 34202 9168 36858
rect 9312 36780 9364 36786
rect 9312 36722 9364 36728
rect 9220 35624 9272 35630
rect 9220 35566 9272 35572
rect 9232 35222 9260 35566
rect 9220 35216 9272 35222
rect 9220 35158 9272 35164
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9232 34082 9260 35158
rect 9140 34054 9260 34082
rect 9034 31920 9090 31929
rect 9034 31855 9090 31864
rect 9140 31822 9168 34054
rect 9324 33114 9352 36722
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9496 36644 9548 36650
rect 9496 36586 9548 36592
rect 9508 33658 9536 36586
rect 9600 35834 9628 36654
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9588 35828 9640 35834
rect 9588 35770 9640 35776
rect 9600 35154 9628 35770
rect 9692 35766 9720 35974
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9588 35148 9640 35154
rect 9588 35090 9640 35096
rect 9588 34944 9640 34950
rect 9588 34886 9640 34892
rect 9496 33652 9548 33658
rect 9496 33594 9548 33600
rect 9404 33448 9456 33454
rect 9404 33390 9456 33396
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9416 32978 9444 33390
rect 9404 32972 9456 32978
rect 9404 32914 9456 32920
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 8944 31816 8996 31822
rect 8944 31758 8996 31764
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 8956 29850 8984 31758
rect 9140 30802 9168 31758
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 9140 30410 9168 30738
rect 9048 30394 9168 30410
rect 9036 30388 9168 30394
rect 9088 30382 9168 30388
rect 9036 30330 9088 30336
rect 8944 29844 8996 29850
rect 8944 29786 8996 29792
rect 8852 29572 8904 29578
rect 8852 29514 8904 29520
rect 8668 29232 8720 29238
rect 8668 29174 8720 29180
rect 8576 28620 8628 28626
rect 8576 28562 8628 28568
rect 8588 27962 8616 28562
rect 8680 28558 8708 29174
rect 9324 28762 9352 32710
rect 9416 32026 9444 32914
rect 9508 32502 9536 33594
rect 9600 33114 9628 34886
rect 9876 33658 9904 37130
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9968 35086 9996 36518
rect 10060 35290 10088 38898
rect 10152 37754 10180 42502
rect 10244 37874 10272 42758
rect 10336 41449 10364 43726
rect 10428 43110 10456 50186
rect 11704 48748 11756 48754
rect 11704 48690 11756 48696
rect 10784 48612 10836 48618
rect 10784 48554 10836 48560
rect 10600 47048 10652 47054
rect 10600 46990 10652 46996
rect 10508 43716 10560 43722
rect 10508 43658 10560 43664
rect 10416 43104 10468 43110
rect 10416 43046 10468 43052
rect 10322 41440 10378 41449
rect 10322 41375 10378 41384
rect 10324 38412 10376 38418
rect 10324 38354 10376 38360
rect 10336 38010 10364 38354
rect 10324 38004 10376 38010
rect 10324 37946 10376 37952
rect 10232 37868 10284 37874
rect 10232 37810 10284 37816
rect 10152 37726 10272 37754
rect 10244 37126 10272 37726
rect 10428 37330 10456 43046
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10416 37324 10468 37330
rect 10416 37266 10468 37272
rect 10140 37120 10192 37126
rect 10140 37062 10192 37068
rect 10232 37120 10284 37126
rect 10232 37062 10284 37068
rect 10152 36922 10180 37062
rect 10140 36916 10192 36922
rect 10140 36858 10192 36864
rect 10232 36712 10284 36718
rect 10232 36654 10284 36660
rect 10140 35760 10192 35766
rect 10140 35702 10192 35708
rect 10048 35284 10100 35290
rect 10048 35226 10100 35232
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 10152 34950 10180 35702
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 10140 34944 10192 34950
rect 10140 34886 10192 34892
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9496 32496 9548 32502
rect 9496 32438 9548 32444
rect 9772 32224 9824 32230
rect 9772 32166 9824 32172
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9402 31920 9458 31929
rect 9402 31855 9458 31864
rect 9496 31884 9548 31890
rect 9416 30598 9444 31855
rect 9496 31826 9548 31832
rect 9508 31754 9536 31826
rect 9508 31726 9628 31754
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 9416 29646 9444 29990
rect 9404 29640 9456 29646
rect 9404 29582 9456 29588
rect 9600 28762 9628 31726
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9692 29782 9720 30126
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 9784 29714 9812 32166
rect 10060 31482 10088 34886
rect 10244 33658 10272 36654
rect 10336 35018 10364 37266
rect 10324 35012 10376 35018
rect 10324 34954 10376 34960
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 10336 33386 10364 34954
rect 10416 33448 10468 33454
rect 10416 33390 10468 33396
rect 10324 33380 10376 33386
rect 10324 33322 10376 33328
rect 10324 31680 10376 31686
rect 10324 31622 10376 31628
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 10336 30666 10364 31622
rect 10324 30660 10376 30666
rect 10324 30602 10376 30608
rect 10336 30326 10364 30602
rect 10324 30320 10376 30326
rect 10324 30262 10376 30268
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8680 28082 8708 28494
rect 8760 28484 8812 28490
rect 8760 28426 8812 28432
rect 8668 28076 8720 28082
rect 8668 28018 8720 28024
rect 8588 27934 8708 27962
rect 8576 26784 8628 26790
rect 8576 26726 8628 26732
rect 8588 25974 8616 26726
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 8484 24132 8536 24138
rect 8484 24074 8536 24080
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7484 22098 7512 22170
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7300 21690 7328 21830
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7208 21542 7420 21570
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 7024 18970 7052 19994
rect 7208 19922 7236 21422
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6932 17678 6960 18158
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 16946 6960 17614
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7300 17270 7328 17546
rect 7288 17264 7340 17270
rect 7288 17206 7340 17212
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6748 16918 6960 16946
rect 6748 15570 6776 16918
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6748 15314 6776 15506
rect 6932 15434 6960 16390
rect 7024 16250 7052 17138
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7300 16046 7328 17206
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6748 15286 6868 15314
rect 6840 13326 6868 15286
rect 6932 15026 6960 15370
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6932 14464 6960 14962
rect 6932 14436 7052 14464
rect 7024 14362 7052 14436
rect 7024 14346 7236 14362
rect 7024 14340 7248 14346
rect 7024 14334 7196 14340
rect 7196 14282 7248 14288
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 8634 6868 13262
rect 7116 9518 7144 13330
rect 7392 12434 7420 21542
rect 7576 21418 7604 22102
rect 7668 21690 7696 22578
rect 7852 22574 7880 23122
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7484 16250 7512 19450
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7576 15162 7604 19314
rect 7668 16658 7696 20810
rect 7760 20602 7788 21830
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7852 20482 7880 22510
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8128 21146 8156 21490
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8312 21010 8340 22918
rect 8404 21706 8432 24006
rect 8496 23610 8524 24074
rect 8496 23582 8616 23610
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8496 21962 8524 23462
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8404 21678 8524 21706
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7852 20466 8064 20482
rect 7748 20460 7800 20466
rect 7852 20460 8076 20466
rect 7852 20454 8024 20460
rect 7748 20402 7800 20408
rect 8024 20402 8076 20408
rect 7760 18834 7788 20402
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 7944 19802 7972 20334
rect 7852 19774 7972 19802
rect 7852 19446 7880 19774
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7852 18630 7880 19382
rect 8496 19378 8524 21678
rect 8588 20806 8616 23582
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8576 20324 8628 20330
rect 8576 20266 8628 20272
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7852 17066 7880 18022
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7840 17060 7892 17066
rect 7760 17020 7840 17048
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 15706 7696 15982
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 13258 7604 14282
rect 7760 13394 7788 17020
rect 7840 17002 7892 17008
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15094 7880 15846
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7300 12406 7420 12434
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6656 6886 6776 6914
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5920 800 5948 2994
rect 6288 800 6316 3470
rect 6472 2650 6500 4762
rect 6748 3738 6776 6886
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6656 800 6684 2382
rect 7024 800 7052 2926
rect 7300 2922 7328 12406
rect 7576 8838 7604 13194
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 8496 5710 8524 19314
rect 8588 18970 8616 20266
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8588 16250 8616 16526
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8588 14278 8616 14894
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8588 14006 8616 14214
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8484 5704 8536 5710
rect 7838 5672 7894 5681
rect 8484 5646 8536 5652
rect 7838 5607 7894 5616
rect 7654 4176 7710 4185
rect 7654 4111 7710 4120
rect 7668 3738 7696 4111
rect 7852 4010 7880 5607
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 8390 3768 8446 3777
rect 7656 3732 7708 3738
rect 8390 3703 8392 3712
rect 7656 3674 7708 3680
rect 8444 3703 8446 3712
rect 8392 3674 8444 3680
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7392 800 7420 3470
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 800 7788 2246
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 3470
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 2926
rect 8680 2582 8708 27934
rect 8772 24070 8800 28426
rect 9692 28218 9720 29038
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 10046 27296 10102 27305
rect 10046 27231 10102 27240
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8956 26042 8984 26726
rect 9324 26586 9352 26930
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 8944 26036 8996 26042
rect 8944 25978 8996 25984
rect 9416 25770 9444 26930
rect 10060 26518 10088 27231
rect 10048 26512 10100 26518
rect 10048 26454 10100 26460
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 9048 23866 9076 25230
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9404 24676 9456 24682
rect 9404 24618 9456 24624
rect 9416 24274 9444 24618
rect 9508 24410 9536 24822
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9048 22982 9076 23598
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9140 22438 9168 24142
rect 9416 23594 9444 24210
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9508 23662 9536 24074
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9404 23588 9456 23594
rect 9404 23530 9456 23536
rect 9692 23050 9720 24754
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8772 14482 8800 14894
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13938 8800 14418
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8956 4214 8984 22170
rect 9508 22030 9536 22918
rect 9692 22710 9720 22986
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9128 21616 9180 21622
rect 9128 21558 9180 21564
rect 9140 20058 9168 21558
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 15162 9168 16526
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9048 14482 9076 14894
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13326 9076 14214
rect 9232 14074 9260 20742
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8864 800 8892 4082
rect 9048 2378 9076 13262
rect 9324 12986 9352 16934
rect 9416 16046 9444 19246
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15366 9444 15982
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9508 14362 9536 21830
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9692 19514 9720 21286
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 16794 9628 17478
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 14618 9628 16594
rect 9692 15162 9720 18294
rect 9784 16250 9812 25094
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 9876 17066 9904 24754
rect 10152 23304 10180 29650
rect 10336 29238 10364 30262
rect 10428 30122 10456 33390
rect 10520 33318 10548 43658
rect 10612 42566 10640 46990
rect 10692 44872 10744 44878
rect 10692 44814 10744 44820
rect 10704 43790 10732 44814
rect 10796 44742 10824 48554
rect 11612 47048 11664 47054
rect 11612 46990 11664 46996
rect 10876 44804 10928 44810
rect 10876 44746 10928 44752
rect 11060 44804 11112 44810
rect 11060 44746 11112 44752
rect 10784 44736 10836 44742
rect 10784 44678 10836 44684
rect 10692 43784 10744 43790
rect 10692 43726 10744 43732
rect 10704 43450 10732 43726
rect 10692 43444 10744 43450
rect 10692 43386 10744 43392
rect 10600 42560 10652 42566
rect 10600 42502 10652 42508
rect 10600 41608 10652 41614
rect 10600 41550 10652 41556
rect 10612 37806 10640 41550
rect 10600 37800 10652 37806
rect 10600 37742 10652 37748
rect 10692 37800 10744 37806
rect 10692 37742 10744 37748
rect 10508 33312 10560 33318
rect 10508 33254 10560 33260
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10520 31822 10548 32370
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10508 31204 10560 31210
rect 10508 31146 10560 31152
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10416 29776 10468 29782
rect 10416 29718 10468 29724
rect 10324 29232 10376 29238
rect 10324 29174 10376 29180
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10244 26042 10272 28970
rect 10336 28218 10364 29174
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10336 24732 10364 28154
rect 10428 27130 10456 29718
rect 10520 27962 10548 31146
rect 10612 29714 10640 37742
rect 10704 37466 10732 37742
rect 10692 37460 10744 37466
rect 10692 37402 10744 37408
rect 10692 35624 10744 35630
rect 10692 35566 10744 35572
rect 10704 31278 10732 35566
rect 10888 34649 10916 44746
rect 11072 44198 11100 44746
rect 11060 44192 11112 44198
rect 11060 44134 11112 44140
rect 11520 42628 11572 42634
rect 11520 42570 11572 42576
rect 11152 42084 11204 42090
rect 11152 42026 11204 42032
rect 11164 40934 11192 42026
rect 11428 42016 11480 42022
rect 11428 41958 11480 41964
rect 11440 41478 11468 41958
rect 11428 41472 11480 41478
rect 11428 41414 11480 41420
rect 11348 41386 11468 41414
rect 11152 40928 11204 40934
rect 11152 40870 11204 40876
rect 11164 39642 11192 40870
rect 11244 39840 11296 39846
rect 11244 39782 11296 39788
rect 11256 39642 11284 39782
rect 11152 39636 11204 39642
rect 11152 39578 11204 39584
rect 11244 39636 11296 39642
rect 11244 39578 11296 39584
rect 11152 38752 11204 38758
rect 11152 38694 11204 38700
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 11072 37874 11100 38150
rect 11164 38010 11192 38694
rect 11244 38480 11296 38486
rect 11244 38422 11296 38428
rect 11256 38214 11284 38422
rect 11348 38418 11376 41386
rect 11428 40452 11480 40458
rect 11428 40394 11480 40400
rect 11440 40186 11468 40394
rect 11428 40180 11480 40186
rect 11428 40122 11480 40128
rect 11336 38412 11388 38418
rect 11336 38354 11388 38360
rect 11336 38276 11388 38282
rect 11336 38218 11388 38224
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 11348 38010 11376 38218
rect 11152 38004 11204 38010
rect 11152 37946 11204 37952
rect 11336 38004 11388 38010
rect 11336 37946 11388 37952
rect 11060 37868 11112 37874
rect 11060 37810 11112 37816
rect 11060 37664 11112 37670
rect 11060 37606 11112 37612
rect 11072 35630 11100 37606
rect 11336 37120 11388 37126
rect 11336 37062 11388 37068
rect 11060 35624 11112 35630
rect 11060 35566 11112 35572
rect 10874 34640 10930 34649
rect 10874 34575 10930 34584
rect 10888 31754 10916 34575
rect 11060 33380 11112 33386
rect 11060 33322 11112 33328
rect 11072 32026 11100 33322
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 10796 31726 10916 31754
rect 10796 31482 10824 31726
rect 10784 31476 10836 31482
rect 10784 31418 10836 31424
rect 10692 31272 10744 31278
rect 10692 31214 10744 31220
rect 10796 31090 10824 31418
rect 10704 31062 10824 31090
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10520 27934 10640 27962
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10520 26382 10548 27406
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10612 26314 10640 27934
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10612 25770 10640 26250
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10336 24704 10456 24732
rect 10428 24138 10456 24704
rect 10416 24132 10468 24138
rect 10416 24074 10468 24080
rect 10152 23276 10272 23304
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10060 21962 10088 22714
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10060 17610 10088 21898
rect 10152 20330 10180 23122
rect 10244 22234 10272 23276
rect 10600 22432 10652 22438
rect 10600 22374 10652 22380
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10152 17338 10180 19654
rect 10244 19514 10272 21490
rect 10416 21480 10468 21486
rect 10414 21448 10416 21457
rect 10468 21448 10470 21457
rect 10414 21383 10470 21392
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10336 20602 10364 20946
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10336 19310 10364 20538
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10612 18426 10640 22374
rect 10704 21690 10732 31062
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 29646 11008 29990
rect 11256 29714 11284 30874
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 11152 29232 11204 29238
rect 11152 29174 11204 29180
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11072 28218 11100 28902
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10784 28008 10836 28014
rect 10784 27950 10836 27956
rect 10796 27130 10824 27950
rect 10876 27940 10928 27946
rect 10876 27882 10928 27888
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10796 26450 10824 27066
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10888 24954 10916 27882
rect 11072 26586 11100 28154
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 11164 26234 11192 29174
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 11256 26994 11284 28494
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11164 26206 11284 26234
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 11060 24744 11112 24750
rect 10980 24704 11060 24732
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10888 23662 10916 24006
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10888 22574 10916 23598
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10980 22438 11008 24704
rect 11060 24686 11112 24692
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 11256 22094 11284 26206
rect 11348 25294 11376 37062
rect 11440 36174 11468 40122
rect 11532 38554 11560 42570
rect 11624 42362 11652 46990
rect 11716 44538 11744 48690
rect 11900 47258 11928 51954
rect 11992 48890 12020 52430
rect 11980 48884 12032 48890
rect 11980 48826 12032 48832
rect 11888 47252 11940 47258
rect 11888 47194 11940 47200
rect 11796 45484 11848 45490
rect 11796 45426 11848 45432
rect 11704 44532 11756 44538
rect 11704 44474 11756 44480
rect 11808 44305 11836 45426
rect 12348 44736 12400 44742
rect 12348 44678 12400 44684
rect 11980 44396 12032 44402
rect 11980 44338 12032 44344
rect 11794 44296 11850 44305
rect 11794 44231 11850 44240
rect 11796 43784 11848 43790
rect 11796 43726 11848 43732
rect 11808 42702 11836 43726
rect 11796 42696 11848 42702
rect 11796 42638 11848 42644
rect 11612 42356 11664 42362
rect 11612 42298 11664 42304
rect 11808 41698 11836 42638
rect 11888 42220 11940 42226
rect 11888 42162 11940 42168
rect 11716 41682 11836 41698
rect 11704 41676 11836 41682
rect 11756 41670 11836 41676
rect 11704 41618 11756 41624
rect 11612 41064 11664 41070
rect 11612 41006 11664 41012
rect 11624 39846 11652 41006
rect 11808 40458 11836 41670
rect 11796 40452 11848 40458
rect 11796 40394 11848 40400
rect 11704 39908 11756 39914
rect 11704 39850 11756 39856
rect 11612 39840 11664 39846
rect 11612 39782 11664 39788
rect 11624 38826 11652 39782
rect 11716 39574 11744 39850
rect 11704 39568 11756 39574
rect 11704 39510 11756 39516
rect 11900 39098 11928 42162
rect 11992 41274 12020 44338
rect 12360 44334 12388 44678
rect 12544 44538 12572 53382
rect 12728 53174 12756 56200
rect 13096 56114 13124 56200
rect 13188 56114 13216 56222
rect 13096 56086 13216 56114
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12716 53168 12768 53174
rect 12716 53110 12768 53116
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 13372 52494 13400 56222
rect 13450 56200 13506 57000
rect 13818 56200 13874 57000
rect 14186 56200 14242 57000
rect 14554 56200 14610 57000
rect 14922 56200 14978 57000
rect 15290 56200 15346 57000
rect 15658 56200 15714 57000
rect 16026 56200 16082 57000
rect 16394 56200 16450 57000
rect 16762 56200 16818 57000
rect 17130 56200 17186 57000
rect 17498 56200 17554 57000
rect 17866 56200 17922 57000
rect 18234 56200 18290 57000
rect 18602 56200 18658 57000
rect 18970 56200 19026 57000
rect 19338 56200 19394 57000
rect 19706 56200 19762 57000
rect 20074 56200 20130 57000
rect 20442 56200 20498 57000
rect 20810 56200 20866 57000
rect 21178 56200 21234 57000
rect 21546 56200 21602 57000
rect 21914 56200 21970 57000
rect 22282 56200 22338 57000
rect 22650 56200 22706 57000
rect 23018 56200 23074 57000
rect 23124 56222 23336 56250
rect 13464 53106 13492 56200
rect 13832 53582 13860 56200
rect 14200 53582 14228 56200
rect 14568 54194 14596 56200
rect 14936 54262 14964 56200
rect 14924 54256 14976 54262
rect 14924 54198 14976 54204
rect 15304 54194 15332 56200
rect 14556 54188 14608 54194
rect 14556 54130 14608 54136
rect 15292 54188 15344 54194
rect 15292 54130 15344 54136
rect 14832 53984 14884 53990
rect 14830 53952 14832 53961
rect 15568 53984 15620 53990
rect 14884 53952 14886 53961
rect 15568 53926 15620 53932
rect 14830 53887 14886 53896
rect 13820 53576 13872 53582
rect 13820 53518 13872 53524
rect 14188 53576 14240 53582
rect 14188 53518 14240 53524
rect 14464 53440 14516 53446
rect 14464 53382 14516 53388
rect 13452 53100 13504 53106
rect 13452 53042 13504 53048
rect 13728 52896 13780 52902
rect 13728 52838 13780 52844
rect 13452 52624 13504 52630
rect 13452 52566 13504 52572
rect 13360 52488 13412 52494
rect 13360 52430 13412 52436
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13360 46504 13412 46510
rect 13360 46446 13412 46452
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 13372 45422 13400 46446
rect 13360 45416 13412 45422
rect 13360 45358 13412 45364
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12532 44532 12584 44538
rect 12532 44474 12584 44480
rect 12716 44396 12768 44402
rect 12716 44338 12768 44344
rect 12164 44328 12216 44334
rect 12164 44270 12216 44276
rect 12348 44328 12400 44334
rect 12348 44270 12400 44276
rect 12176 43450 12204 44270
rect 12256 44192 12308 44198
rect 12256 44134 12308 44140
rect 12268 43602 12296 44134
rect 12360 43722 12388 44270
rect 12348 43716 12400 43722
rect 12348 43658 12400 43664
rect 12268 43574 12388 43602
rect 12164 43444 12216 43450
rect 12164 43386 12216 43392
rect 12360 43178 12388 43574
rect 12348 43172 12400 43178
rect 12348 43114 12400 43120
rect 12256 42288 12308 42294
rect 12256 42230 12308 42236
rect 12072 41540 12124 41546
rect 12072 41482 12124 41488
rect 12084 41290 12112 41482
rect 12084 41274 12204 41290
rect 11980 41268 12032 41274
rect 11980 41210 12032 41216
rect 12072 41268 12204 41274
rect 12124 41262 12204 41268
rect 12072 41210 12124 41216
rect 12072 41132 12124 41138
rect 12072 41074 12124 41080
rect 11888 39092 11940 39098
rect 11888 39034 11940 39040
rect 11612 38820 11664 38826
rect 11612 38762 11664 38768
rect 11520 38548 11572 38554
rect 11520 38490 11572 38496
rect 11520 37800 11572 37806
rect 11520 37742 11572 37748
rect 11532 37398 11560 37742
rect 12084 37738 12112 41074
rect 12176 40594 12204 41262
rect 12164 40588 12216 40594
rect 12164 40530 12216 40536
rect 12164 40452 12216 40458
rect 12164 40394 12216 40400
rect 12176 39982 12204 40394
rect 12164 39976 12216 39982
rect 12164 39918 12216 39924
rect 12176 39506 12204 39918
rect 12164 39500 12216 39506
rect 12164 39442 12216 39448
rect 12268 39370 12296 42230
rect 12360 41070 12388 43114
rect 12624 42764 12676 42770
rect 12624 42706 12676 42712
rect 12636 41478 12664 42706
rect 12624 41472 12676 41478
rect 12624 41414 12676 41420
rect 12348 41064 12400 41070
rect 12348 41006 12400 41012
rect 12624 40588 12676 40594
rect 12624 40530 12676 40536
rect 12348 40452 12400 40458
rect 12348 40394 12400 40400
rect 12360 40066 12388 40394
rect 12532 40180 12584 40186
rect 12532 40122 12584 40128
rect 12440 40112 12492 40118
rect 12360 40060 12440 40066
rect 12360 40054 12492 40060
rect 12360 40038 12480 40054
rect 12360 39438 12388 40038
rect 12544 39982 12572 40122
rect 12440 39976 12492 39982
rect 12440 39918 12492 39924
rect 12532 39976 12584 39982
rect 12532 39918 12584 39924
rect 12452 39506 12480 39918
rect 12440 39500 12492 39506
rect 12440 39442 12492 39448
rect 12348 39432 12400 39438
rect 12348 39374 12400 39380
rect 12256 39364 12308 39370
rect 12256 39306 12308 39312
rect 12164 39296 12216 39302
rect 12164 39238 12216 39244
rect 12348 39296 12400 39302
rect 12348 39238 12400 39244
rect 12176 38486 12204 39238
rect 12256 38888 12308 38894
rect 12256 38830 12308 38836
rect 12164 38480 12216 38486
rect 12164 38422 12216 38428
rect 12072 37732 12124 37738
rect 12072 37674 12124 37680
rect 12176 37670 12204 38422
rect 12164 37664 12216 37670
rect 12164 37606 12216 37612
rect 11520 37392 11572 37398
rect 11520 37334 11572 37340
rect 11428 36168 11480 36174
rect 11428 36110 11480 36116
rect 11532 31754 11560 37334
rect 11796 36100 11848 36106
rect 11796 36042 11848 36048
rect 11808 35630 11836 36042
rect 11886 36000 11942 36009
rect 11886 35935 11942 35944
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11808 35222 11836 35566
rect 11796 35216 11848 35222
rect 11796 35158 11848 35164
rect 11808 34626 11836 35158
rect 11716 34610 11836 34626
rect 11704 34604 11836 34610
rect 11756 34598 11836 34604
rect 11704 34546 11756 34552
rect 11704 34128 11756 34134
rect 11704 34070 11756 34076
rect 11440 31726 11560 31754
rect 11440 30546 11468 31726
rect 11440 30518 11560 30546
rect 11428 26988 11480 26994
rect 11428 26930 11480 26936
rect 11440 25838 11468 26930
rect 11428 25832 11480 25838
rect 11428 25774 11480 25780
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11532 24698 11560 30518
rect 11716 25158 11744 34070
rect 11900 33930 11928 35935
rect 11992 34870 12204 34898
rect 11992 34746 12020 34870
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 11888 33924 11940 33930
rect 11888 33866 11940 33872
rect 11900 33833 11928 33866
rect 11980 33856 12032 33862
rect 11886 33824 11942 33833
rect 11980 33798 12032 33804
rect 11886 33759 11942 33768
rect 11992 32026 12020 33798
rect 12084 32774 12112 34682
rect 12176 33130 12204 34870
rect 12268 34202 12296 38830
rect 12360 38418 12388 39238
rect 12348 38412 12400 38418
rect 12348 38354 12400 38360
rect 12348 38208 12400 38214
rect 12348 38150 12400 38156
rect 12256 34196 12308 34202
rect 12256 34138 12308 34144
rect 12360 34134 12388 38150
rect 12452 36258 12480 39442
rect 12532 39432 12584 39438
rect 12532 39374 12584 39380
rect 12544 36378 12572 39374
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 12636 36360 12664 40530
rect 12728 39438 12756 44338
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13372 42158 13400 45358
rect 13360 42152 13412 42158
rect 13360 42094 13412 42100
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 13372 41682 13400 42094
rect 13360 41676 13412 41682
rect 13360 41618 13412 41624
rect 13372 41138 13400 41618
rect 13360 41132 13412 41138
rect 13360 41074 13412 41080
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 13464 40526 13492 52566
rect 13636 45552 13688 45558
rect 13636 45494 13688 45500
rect 13544 43648 13596 43654
rect 13544 43590 13596 43596
rect 13452 40520 13504 40526
rect 13452 40462 13504 40468
rect 13556 39914 13584 43590
rect 13544 39908 13596 39914
rect 13544 39850 13596 39856
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 13556 39438 13584 39850
rect 13648 39642 13676 45494
rect 13636 39636 13688 39642
rect 13636 39578 13688 39584
rect 12716 39432 12768 39438
rect 12716 39374 12768 39380
rect 13544 39432 13596 39438
rect 13544 39374 13596 39380
rect 12992 39296 13044 39302
rect 12992 39238 13044 39244
rect 13004 39030 13032 39238
rect 12716 39024 12768 39030
rect 12716 38966 12768 38972
rect 12992 39024 13044 39030
rect 12992 38966 13044 38972
rect 12728 36922 12756 38966
rect 13360 38752 13412 38758
rect 13360 38694 13412 38700
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 13372 38418 13400 38694
rect 13360 38412 13412 38418
rect 13360 38354 13412 38360
rect 12808 38004 12860 38010
rect 12808 37946 12860 37952
rect 12820 37670 12848 37946
rect 12808 37664 12860 37670
rect 12808 37606 12860 37612
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13084 36372 13136 36378
rect 12636 36332 12848 36360
rect 12452 36230 12572 36258
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12348 34128 12400 34134
rect 12348 34070 12400 34076
rect 12256 34060 12308 34066
rect 12256 34002 12308 34008
rect 12268 33862 12296 34002
rect 12348 33992 12400 33998
rect 12452 33980 12480 35974
rect 12544 34066 12572 36230
rect 12636 34542 12664 36332
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12624 34536 12676 34542
rect 12624 34478 12676 34484
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12400 33952 12480 33980
rect 12348 33934 12400 33940
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 12624 33312 12676 33318
rect 12624 33254 12676 33260
rect 12176 33102 12296 33130
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 12072 32768 12124 32774
rect 12072 32710 12124 32716
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 12176 29782 12204 32846
rect 12268 30870 12296 33102
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 12164 29776 12216 29782
rect 12164 29718 12216 29724
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 11888 28144 11940 28150
rect 11888 28086 11940 28092
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 11704 25152 11756 25158
rect 11704 25094 11756 25100
rect 11532 24670 11652 24698
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11256 22066 11376 22094
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10704 20806 10732 21626
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10980 18970 11008 21422
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 19514 11100 20266
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11164 19854 11192 20198
rect 11256 19922 11284 20198
rect 11348 19922 11376 22066
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10980 18442 11008 18906
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10796 18414 11008 18442
rect 11072 18426 11100 19450
rect 11060 18420 11112 18426
rect 10796 18272 10824 18414
rect 11060 18362 11112 18368
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10520 18244 10824 18272
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10244 17610 10272 18022
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 10244 16794 10272 17546
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 9772 16244 9824 16250
rect 9824 16204 9904 16232
rect 9772 16186 9824 16192
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9416 12238 9444 14350
rect 9508 14334 9720 14362
rect 9692 14278 9720 14334
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11694 9444 12174
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9232 800 9260 4082
rect 9416 3058 9444 4966
rect 9508 4010 9536 14010
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12782 9720 13126
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12306 9720 12718
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9600 3738 9628 5510
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9508 2514 9536 2790
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 800 9628 3470
rect 9784 2446 9812 14894
rect 9876 10062 9904 16204
rect 10244 15502 10272 16730
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 16046 10364 16594
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10048 15156 10100 15162
rect 10100 15116 10180 15144
rect 10048 15098 10100 15104
rect 10152 14006 10180 15116
rect 10244 14414 10272 15438
rect 10336 14822 10364 15982
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10336 14346 10364 14758
rect 10520 14618 10548 18244
rect 10888 18170 10916 18294
rect 10612 18142 10916 18170
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10152 12170 10180 13942
rect 10520 13938 10548 14554
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 11082 10180 12106
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 10612 6914 10640 18142
rect 11072 17134 11100 18362
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11164 16674 11192 19654
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18834 11376 19110
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10888 16646 11192 16674
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16182 10732 16390
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10796 14006 10824 16594
rect 10888 16590 10916 16646
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16250 10916 16390
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11072 15434 11100 16458
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 15162 11100 15370
rect 11060 15156 11112 15162
rect 11112 15116 11192 15144
rect 11060 15098 11112 15104
rect 11164 14346 11192 15116
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10336 6886 10640 6914
rect 10336 5574 10364 6886
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9968 800 9996 3470
rect 10612 3058 10640 5578
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 10336 800 10364 2926
rect 10704 800 10732 3470
rect 10796 2650 10824 13942
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10888 11286 10916 13874
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12306 11008 12582
rect 11164 12442 11192 13330
rect 11152 12436 11204 12442
rect 11256 12434 11284 18566
rect 11348 18222 11376 18770
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11348 16590 11376 16730
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 11440 14822 11468 22918
rect 11532 20942 11560 24006
rect 11624 23798 11652 24670
rect 11612 23792 11664 23798
rect 11612 23734 11664 23740
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11624 20890 11652 22102
rect 11716 21554 11744 25094
rect 11808 22574 11836 25774
rect 11900 23610 11928 28086
rect 12070 27976 12126 27985
rect 12070 27911 12126 27920
rect 12084 27062 12112 27911
rect 12176 27418 12204 29582
rect 12360 28218 12388 32166
rect 12636 30598 12664 33254
rect 12728 33046 12756 36178
rect 12820 35834 12848 36332
rect 13084 36314 13136 36320
rect 12808 35828 12860 35834
rect 12808 35770 12860 35776
rect 13096 35562 13124 36314
rect 13372 36174 13400 38354
rect 13636 37256 13688 37262
rect 13636 37198 13688 37204
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 13452 36712 13504 36718
rect 13452 36654 13504 36660
rect 13360 36168 13412 36174
rect 13360 36110 13412 36116
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 13084 35556 13136 35562
rect 13084 35498 13136 35504
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 13372 35086 13400 35634
rect 13464 35494 13492 36654
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13452 35216 13504 35222
rect 13452 35158 13504 35164
rect 13360 35080 13412 35086
rect 13360 35022 13412 35028
rect 13372 34678 13400 35022
rect 13360 34672 13412 34678
rect 13360 34614 13412 34620
rect 13360 34536 13412 34542
rect 13360 34478 13412 34484
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 13268 33924 13320 33930
rect 13268 33866 13320 33872
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 12820 33658 12848 33798
rect 12808 33652 12860 33658
rect 12808 33594 12860 33600
rect 13280 33318 13308 33866
rect 13372 33386 13400 34478
rect 13464 34066 13492 35158
rect 13452 34060 13504 34066
rect 13452 34002 13504 34008
rect 13360 33380 13412 33386
rect 13360 33322 13412 33328
rect 13268 33312 13320 33318
rect 13268 33254 13320 33260
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12716 33040 12768 33046
rect 12716 32982 12768 32988
rect 12728 31890 12756 32982
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13280 32434 13308 32710
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12716 31680 12768 31686
rect 12714 31648 12716 31657
rect 12768 31648 12770 31657
rect 12714 31583 12770 31592
rect 12532 30592 12584 30598
rect 12532 30534 12584 30540
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12452 29306 12480 29650
rect 12544 29578 12572 30534
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12532 29572 12584 29578
rect 12532 29514 12584 29520
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 12348 27872 12400 27878
rect 12348 27814 12400 27820
rect 12254 27432 12310 27441
rect 12176 27390 12254 27418
rect 12254 27367 12310 27376
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11992 24426 12020 26726
rect 12070 24984 12126 24993
rect 12070 24919 12072 24928
rect 12124 24919 12126 24928
rect 12072 24890 12124 24896
rect 11992 24398 12112 24426
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 23798 12020 24006
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11900 23594 12020 23610
rect 11900 23588 12032 23594
rect 11900 23582 11980 23588
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11808 22098 11836 22510
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11624 20862 11744 20890
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11624 19514 11652 20742
rect 11716 19718 11744 20862
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11532 15706 11560 17818
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11256 12406 11376 12434
rect 11152 12378 11204 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 11164 11082 11192 12378
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11218 11284 11630
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11348 6914 11376 12406
rect 11256 6886 11376 6914
rect 11256 6254 11284 6886
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11624 4826 11652 18770
rect 11716 18426 11744 19314
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 12986 11744 17138
rect 11808 14618 11836 19382
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11900 12238 11928 23582
rect 11980 23530 12032 23536
rect 12084 22506 12112 24398
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12176 22522 12204 24210
rect 12268 22982 12296 27367
rect 12360 23866 12388 27814
rect 12452 25265 12480 28970
rect 12544 28626 12572 29514
rect 12636 29034 12664 29786
rect 12624 29028 12676 29034
rect 12624 28970 12676 28976
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 12636 28082 12664 28494
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12636 27674 12664 28018
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12532 27600 12584 27606
rect 12532 27542 12584 27548
rect 12438 25256 12494 25265
rect 12438 25191 12494 25200
rect 12440 24948 12492 24954
rect 12544 24936 12572 27542
rect 12544 24908 12664 24936
rect 12440 24890 12492 24896
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12072 22500 12124 22506
rect 12176 22494 12296 22522
rect 12072 22442 12124 22448
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11992 21146 12020 21422
rect 12084 21418 12112 21927
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 12084 21010 12112 21354
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12176 20602 12204 22374
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12268 20482 12296 22494
rect 12348 21888 12400 21894
rect 12346 21856 12348 21865
rect 12400 21856 12402 21865
rect 12346 21791 12402 21800
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12084 20454 12296 20482
rect 12084 20398 12112 20454
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11992 17746 12020 19858
rect 12084 19446 12112 20334
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12084 17338 12112 18566
rect 12176 18154 12204 20334
rect 12360 20058 12388 21490
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12268 16658 12296 19654
rect 12452 19530 12480 24890
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12360 19502 12480 19530
rect 12360 18698 12388 19502
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12544 18578 12572 24754
rect 12636 22710 12664 24908
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12728 22094 12756 31583
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 13372 30938 13400 33322
rect 13556 33318 13584 36722
rect 13648 35834 13676 37198
rect 13636 35828 13688 35834
rect 13636 35770 13688 35776
rect 13634 35184 13690 35193
rect 13634 35119 13636 35128
rect 13688 35119 13690 35128
rect 13636 35090 13688 35096
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13544 33312 13596 33318
rect 13544 33254 13596 33260
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 13360 30592 13412 30598
rect 13358 30560 13360 30569
rect 13412 30560 13414 30569
rect 13358 30495 13414 30504
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 13004 30161 13032 30194
rect 12990 30152 13046 30161
rect 12990 30087 13046 30096
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13372 29850 13400 30330
rect 13360 29844 13412 29850
rect 13360 29786 13412 29792
rect 13464 29714 13492 33254
rect 13648 32910 13676 35090
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12912 29034 12940 29446
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 12900 29028 12952 29034
rect 12900 28970 12952 28976
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 12820 26874 12848 28358
rect 13372 28150 13400 29242
rect 13360 28144 13412 28150
rect 13360 28086 13412 28092
rect 13360 27872 13412 27878
rect 13360 27814 13412 27820
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 13096 26994 13124 27610
rect 13176 27464 13228 27470
rect 13372 27452 13400 27814
rect 13228 27424 13400 27452
rect 13176 27406 13228 27412
rect 13176 27328 13228 27334
rect 13174 27296 13176 27305
rect 13228 27296 13230 27305
rect 13230 27254 13400 27282
rect 13174 27231 13230 27240
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12820 26858 13032 26874
rect 12820 26852 13044 26858
rect 12820 26846 12992 26852
rect 12820 25838 12848 26846
rect 12992 26794 13044 26800
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13188 25906 13216 26522
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12820 25362 12848 25774
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12806 25256 12862 25265
rect 12806 25191 12862 25200
rect 12820 22658 12848 25191
rect 12898 25120 12954 25129
rect 12898 25055 12954 25064
rect 12912 24818 12940 25055
rect 13372 24818 13400 27254
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13464 26234 13492 26862
rect 13556 26382 13584 29990
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13464 26206 13584 26234
rect 13556 25702 13584 26206
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13556 24342 13584 25638
rect 13648 24954 13676 32846
rect 13740 29306 13768 52838
rect 14096 52488 14148 52494
rect 14096 52430 14148 52436
rect 13820 44736 13872 44742
rect 13820 44678 13872 44684
rect 13832 43790 13860 44678
rect 13820 43784 13872 43790
rect 13820 43726 13872 43732
rect 13820 42900 13872 42906
rect 13820 42842 13872 42848
rect 13832 41052 13860 42842
rect 13912 42016 13964 42022
rect 13912 41958 13964 41964
rect 13924 41206 13952 41958
rect 13912 41200 13964 41206
rect 13912 41142 13964 41148
rect 14004 41064 14056 41070
rect 13832 41024 14004 41052
rect 13832 40746 13860 41024
rect 14004 41006 14056 41012
rect 13832 40718 13952 40746
rect 13820 40656 13872 40662
rect 13820 40598 13872 40604
rect 13832 38978 13860 40598
rect 13924 40118 13952 40718
rect 13912 40112 13964 40118
rect 13912 40054 13964 40060
rect 13912 39840 13964 39846
rect 13912 39782 13964 39788
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 13924 39506 13952 39782
rect 13912 39500 13964 39506
rect 13912 39442 13964 39448
rect 14016 39098 14044 39782
rect 14004 39092 14056 39098
rect 14004 39034 14056 39040
rect 13832 38950 13952 38978
rect 13820 38888 13872 38894
rect 13820 38830 13872 38836
rect 13832 37738 13860 38830
rect 13820 37732 13872 37738
rect 13820 37674 13872 37680
rect 13820 35080 13872 35086
rect 13820 35022 13872 35028
rect 13832 32978 13860 35022
rect 13924 33658 13952 38950
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 14016 33862 14044 35430
rect 14004 33856 14056 33862
rect 14004 33798 14056 33804
rect 13912 33652 13964 33658
rect 13912 33594 13964 33600
rect 14004 33584 14056 33590
rect 14004 33526 14056 33532
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 14016 31754 14044 33526
rect 13832 31726 14044 31754
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13728 26512 13780 26518
rect 13728 26454 13780 26460
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13096 23866 13124 24074
rect 13464 23866 13492 24142
rect 13648 23866 13676 24754
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12820 22642 12940 22658
rect 12820 22636 12952 22642
rect 12820 22630 12900 22636
rect 12900 22578 12952 22584
rect 12808 22568 12860 22574
rect 12912 22545 12940 22578
rect 13360 22568 13412 22574
rect 12808 22510 12860 22516
rect 12898 22536 12954 22545
rect 12820 22216 12848 22510
rect 13360 22510 13412 22516
rect 12898 22471 12954 22480
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12820 22188 12940 22216
rect 12728 22066 12848 22094
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12636 21078 12664 21966
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12452 18550 12572 18578
rect 12346 18456 12402 18465
rect 12346 18391 12402 18400
rect 12360 18358 12388 18391
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12360 15978 12388 17070
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11992 12050 12020 13874
rect 11900 12022 12020 12050
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11532 3738 11560 4150
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11072 800 11100 2790
rect 11716 2514 11744 9862
rect 11900 6914 11928 12022
rect 11980 11620 12032 11626
rect 11980 11562 12032 11568
rect 11992 11082 12020 11562
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11900 6886 12020 6914
rect 11992 3058 12020 6886
rect 12084 6390 12112 15642
rect 12360 14278 12388 15914
rect 12452 15094 12480 18550
rect 12636 18222 12664 19246
rect 12728 18766 12756 21830
rect 12820 18834 12848 22066
rect 12912 21554 12940 22188
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 21622 13308 21830
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21010 13400 22510
rect 13556 21978 13584 23666
rect 13740 23050 13768 26454
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13648 22098 13676 22646
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13556 21950 13676 21978
rect 13452 21480 13504 21486
rect 13450 21448 13452 21457
rect 13504 21448 13506 21457
rect 13450 21383 13506 21392
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12912 19174 12940 19994
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 16454 12572 17478
rect 12636 16794 12664 18158
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 12782 12388 14214
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12452 12434 12480 14826
rect 12636 14550 12664 16730
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12728 14074 12756 17002
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15162 12848 16050
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13372 15688 13400 19790
rect 13464 18834 13492 20334
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13556 18698 13584 19314
rect 13544 18692 13596 18698
rect 13544 18634 13596 18640
rect 13556 18578 13584 18634
rect 13280 15660 13400 15688
rect 13464 18550 13584 18578
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12820 14482 12848 14894
rect 13280 14890 13308 15660
rect 13464 15586 13492 18550
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13556 18086 13584 18362
rect 13648 18272 13676 21950
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13740 21146 13768 21490
rect 13832 21468 13860 31726
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 13924 22030 13952 27270
rect 14016 27130 14044 30058
rect 14108 29850 14136 52430
rect 14280 44872 14332 44878
rect 14280 44814 14332 44820
rect 14188 44192 14240 44198
rect 14188 44134 14240 44140
rect 14200 37942 14228 44134
rect 14292 42770 14320 44814
rect 14280 42764 14332 42770
rect 14280 42706 14332 42712
rect 14280 42628 14332 42634
rect 14280 42570 14332 42576
rect 14292 42276 14320 42570
rect 14372 42288 14424 42294
rect 14292 42248 14372 42276
rect 14372 42230 14424 42236
rect 14384 41478 14412 42230
rect 14372 41472 14424 41478
rect 14372 41414 14424 41420
rect 14292 41386 14412 41414
rect 14292 41206 14320 41386
rect 14280 41200 14332 41206
rect 14280 41142 14332 41148
rect 14292 40458 14320 41142
rect 14280 40452 14332 40458
rect 14280 40394 14332 40400
rect 14280 40112 14332 40118
rect 14280 40054 14332 40060
rect 14188 37936 14240 37942
rect 14188 37878 14240 37884
rect 14188 37800 14240 37806
rect 14292 37754 14320 40054
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14240 37748 14320 37754
rect 14188 37742 14320 37748
rect 14200 37726 14320 37742
rect 14384 36922 14412 38150
rect 14372 36916 14424 36922
rect 14372 36858 14424 36864
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14200 34950 14228 35566
rect 14188 34944 14240 34950
rect 14188 34886 14240 34892
rect 14200 33454 14228 34886
rect 14476 34762 14504 53382
rect 14556 52964 14608 52970
rect 14556 52906 14608 52912
rect 14568 52601 14596 52906
rect 14554 52592 14610 52601
rect 14554 52527 14610 52536
rect 15016 46912 15068 46918
rect 15016 46854 15068 46860
rect 15028 46578 15056 46854
rect 15384 46708 15436 46714
rect 15384 46650 15436 46656
rect 15016 46572 15068 46578
rect 15016 46514 15068 46520
rect 15028 45558 15056 46514
rect 15016 45552 15068 45558
rect 15016 45494 15068 45500
rect 15028 44810 15056 45494
rect 15396 45422 15424 46650
rect 15580 46073 15608 53926
rect 15672 53582 15700 56200
rect 16040 54262 16068 56200
rect 16028 54256 16080 54262
rect 16028 54198 16080 54204
rect 15752 54052 15804 54058
rect 15752 53994 15804 54000
rect 15660 53576 15712 53582
rect 15660 53518 15712 53524
rect 15764 51074 15792 53994
rect 16120 53984 16172 53990
rect 16120 53926 16172 53932
rect 15936 53440 15988 53446
rect 15936 53382 15988 53388
rect 15672 51046 15792 51074
rect 15566 46064 15622 46073
rect 15566 45999 15622 46008
rect 15384 45416 15436 45422
rect 15384 45358 15436 45364
rect 15108 45280 15160 45286
rect 15108 45222 15160 45228
rect 14556 44804 14608 44810
rect 14556 44746 14608 44752
rect 15016 44804 15068 44810
rect 15016 44746 15068 44752
rect 14568 44198 14596 44746
rect 14924 44328 14976 44334
rect 14924 44270 14976 44276
rect 14556 44192 14608 44198
rect 14556 44134 14608 44140
rect 14568 38894 14596 44134
rect 14936 42022 14964 44270
rect 15120 42906 15148 45222
rect 15476 44532 15528 44538
rect 15476 44474 15528 44480
rect 15292 43784 15344 43790
rect 15292 43726 15344 43732
rect 15200 43308 15252 43314
rect 15200 43250 15252 43256
rect 15108 42900 15160 42906
rect 15108 42842 15160 42848
rect 14924 42016 14976 42022
rect 14924 41958 14976 41964
rect 15108 41268 15160 41274
rect 15108 41210 15160 41216
rect 14924 40928 14976 40934
rect 14924 40870 14976 40876
rect 14556 38888 14608 38894
rect 14556 38830 14608 38836
rect 14556 38344 14608 38350
rect 14556 38286 14608 38292
rect 14384 34734 14504 34762
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 14292 32065 14320 32166
rect 14278 32056 14334 32065
rect 14278 31991 14334 32000
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14096 29844 14148 29850
rect 14096 29786 14148 29792
rect 14108 28082 14136 29786
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14004 27124 14056 27130
rect 14004 27066 14056 27072
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14016 26586 14044 26930
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13912 21616 13964 21622
rect 13910 21584 13912 21593
rect 13964 21584 13966 21593
rect 13910 21519 13966 21528
rect 13832 21440 14044 21468
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20602 13860 21286
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13728 18284 13780 18290
rect 13648 18244 13728 18272
rect 13728 18226 13780 18232
rect 13544 18080 13596 18086
rect 13596 18040 13676 18068
rect 13544 18022 13596 18028
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 16454 13584 17682
rect 13648 17338 13676 18040
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13740 17134 13768 18226
rect 13924 17270 13952 21286
rect 13912 17264 13964 17270
rect 13912 17206 13964 17212
rect 13728 17128 13780 17134
rect 14016 17082 14044 21440
rect 13728 17070 13780 17076
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13372 15558 13492 15586
rect 13372 15026 13400 15558
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12452 12406 12664 12434
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 12452 3058 12480 12038
rect 12636 5030 12664 12406
rect 12728 8566 12756 13806
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12820 11082 12848 12854
rect 13280 12764 13308 13466
rect 13372 12918 13400 14758
rect 13464 14346 13492 14962
rect 13556 14958 13584 16390
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13464 14074 13492 14282
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13938 13492 14010
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13556 13530 13584 14758
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13280 12736 13400 12764
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12170 13400 12736
rect 13464 12374 13492 13398
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13556 11286 13584 12786
rect 13648 12442 13676 15030
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 12808 11076 12860 11082
rect 12808 11018 12860 11024
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13648 4146 13676 12174
rect 13740 4214 13768 17070
rect 13832 17054 14044 17082
rect 13832 13326 13860 17054
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 14414 13952 16934
rect 14002 16280 14058 16289
rect 14002 16215 14058 16224
rect 14016 16182 14044 16215
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 14108 14958 14136 26930
rect 14200 26450 14228 30534
rect 14292 28626 14320 30670
rect 14384 30258 14412 34734
rect 14568 34406 14596 38286
rect 14936 37806 14964 40870
rect 15016 39976 15068 39982
rect 15016 39918 15068 39924
rect 14924 37800 14976 37806
rect 14844 37748 14924 37754
rect 14844 37742 14976 37748
rect 14844 37726 14964 37742
rect 14648 35488 14700 35494
rect 14648 35430 14700 35436
rect 14556 34400 14608 34406
rect 14556 34342 14608 34348
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14476 31890 14504 32302
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14464 31884 14516 31890
rect 14464 31826 14516 31832
rect 14568 31754 14596 32166
rect 14476 31726 14596 31754
rect 14476 30666 14504 31726
rect 14464 30660 14516 30666
rect 14464 30602 14516 30608
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14384 29238 14412 30194
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14188 26444 14240 26450
rect 14188 26386 14240 26392
rect 14292 24562 14320 28018
rect 14372 27940 14424 27946
rect 14372 27882 14424 27888
rect 14384 24682 14412 27882
rect 14476 27538 14504 30602
rect 14660 30190 14688 35430
rect 14844 35086 14872 37726
rect 14924 37664 14976 37670
rect 14924 37606 14976 37612
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 14832 34468 14884 34474
rect 14832 34410 14884 34416
rect 14740 34128 14792 34134
rect 14740 34070 14792 34076
rect 14752 33590 14780 34070
rect 14740 33584 14792 33590
rect 14740 33526 14792 33532
rect 14740 32768 14792 32774
rect 14740 32710 14792 32716
rect 14648 30184 14700 30190
rect 14648 30126 14700 30132
rect 14556 29164 14608 29170
rect 14556 29106 14608 29112
rect 14464 27532 14516 27538
rect 14464 27474 14516 27480
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14476 25294 14504 26318
rect 14568 25770 14596 29106
rect 14752 27538 14780 32710
rect 14844 32570 14872 34410
rect 14936 33658 14964 37606
rect 15028 34678 15056 39918
rect 15120 35834 15148 41210
rect 15212 40730 15240 43250
rect 15304 42226 15332 43726
rect 15384 43104 15436 43110
rect 15384 43046 15436 43052
rect 15292 42220 15344 42226
rect 15292 42162 15344 42168
rect 15304 41682 15332 42162
rect 15292 41676 15344 41682
rect 15292 41618 15344 41624
rect 15200 40724 15252 40730
rect 15200 40666 15252 40672
rect 15200 39840 15252 39846
rect 15200 39782 15252 39788
rect 15212 39438 15240 39782
rect 15200 39432 15252 39438
rect 15200 39374 15252 39380
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15304 37777 15332 37810
rect 15290 37768 15346 37777
rect 15290 37703 15346 37712
rect 15396 37398 15424 43046
rect 15384 37392 15436 37398
rect 15384 37334 15436 37340
rect 15292 37188 15344 37194
rect 15292 37130 15344 37136
rect 15304 36922 15332 37130
rect 15488 37126 15516 44474
rect 15672 41414 15700 51046
rect 15752 47116 15804 47122
rect 15752 47058 15804 47064
rect 15764 46866 15792 47058
rect 15764 46838 15884 46866
rect 15856 45966 15884 46838
rect 15844 45960 15896 45966
rect 15844 45902 15896 45908
rect 15856 45626 15884 45902
rect 15844 45620 15896 45626
rect 15844 45562 15896 45568
rect 15856 43790 15884 45562
rect 15844 43784 15896 43790
rect 15844 43726 15896 43732
rect 15672 41386 15792 41414
rect 15764 40390 15792 41386
rect 15752 40384 15804 40390
rect 15752 40326 15804 40332
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15292 36916 15344 36922
rect 15292 36858 15344 36864
rect 15290 36272 15346 36281
rect 15290 36207 15346 36216
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 15108 35828 15160 35834
rect 15108 35770 15160 35776
rect 15212 35086 15240 36110
rect 15304 36038 15332 36207
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 15120 33522 15148 34342
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 15028 33114 15056 33458
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 15016 33108 15068 33114
rect 15016 33050 15068 33056
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14844 29646 14872 32506
rect 15016 30320 15068 30326
rect 15016 30262 15068 30268
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14936 29850 14964 29990
rect 14924 29844 14976 29850
rect 14924 29786 14976 29792
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14936 27554 14964 28970
rect 15028 27690 15056 30262
rect 15120 27946 15148 33254
rect 15304 31754 15332 35566
rect 15292 31748 15344 31754
rect 15292 31690 15344 31696
rect 15384 31748 15436 31754
rect 15384 31690 15436 31696
rect 15200 31680 15252 31686
rect 15200 31622 15252 31628
rect 15212 30666 15240 31622
rect 15304 31278 15332 31690
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15212 28506 15240 30602
rect 15292 30184 15344 30190
rect 15290 30152 15292 30161
rect 15344 30152 15346 30161
rect 15290 30087 15346 30096
rect 15396 28762 15424 31690
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15212 28490 15424 28506
rect 15212 28484 15436 28490
rect 15212 28478 15384 28484
rect 15384 28426 15436 28432
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15028 27674 15332 27690
rect 15028 27668 15344 27674
rect 15028 27662 15292 27668
rect 15292 27610 15344 27616
rect 14740 27532 14792 27538
rect 14936 27526 15240 27554
rect 14740 27474 14792 27480
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15120 26926 15148 27066
rect 15108 26920 15160 26926
rect 15106 26888 15108 26897
rect 15160 26888 15162 26897
rect 15106 26823 15162 26832
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14476 24818 14504 25230
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14292 24534 14412 24562
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14200 20942 14228 23802
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 14108 13938 14136 14894
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 11354 13860 11834
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14200 9654 14228 18702
rect 14292 17678 14320 22102
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 15348 14320 17070
rect 14384 15502 14412 24534
rect 14568 24070 14596 25366
rect 14660 24274 14688 26726
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15212 25922 15240 27526
rect 15304 26042 15332 27610
rect 15396 26586 15424 28426
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22778 14504 22918
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 14464 21480 14516 21486
rect 14568 21457 14596 22714
rect 14660 21950 14872 21978
rect 14660 21894 14688 21950
rect 14844 21894 14872 21950
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14752 21690 14780 21830
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14464 21422 14516 21428
rect 14554 21448 14610 21457
rect 14476 20398 14504 21422
rect 14554 21383 14610 21392
rect 14568 21010 14596 21383
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18222 14504 19110
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17134 14504 18158
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 17338 14688 17478
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14752 17270 14780 20198
rect 14844 19700 14872 21830
rect 14936 21554 14964 25638
rect 15120 25498 15148 25910
rect 15212 25894 15424 25922
rect 15108 25492 15160 25498
rect 15108 25434 15160 25440
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15028 20992 15056 24550
rect 14936 20964 15056 20992
rect 14936 19854 14964 20964
rect 15120 20602 15148 25094
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21690 15240 21966
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14844 19672 14964 19700
rect 14740 17264 14792 17270
rect 14740 17206 14792 17212
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14464 15360 14516 15366
rect 14292 15320 14412 15348
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 12850 14320 14418
rect 14384 13802 14412 15320
rect 14464 15302 14516 15308
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11440 800 11468 2382
rect 11808 800 11836 2926
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12176 800 12204 2314
rect 12544 800 12572 3538
rect 12820 2122 12848 4014
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 2094 12940 2122
rect 12912 800 12940 2094
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 14016 800 14044 3538
rect 14292 3534 14320 12650
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14384 11286 14412 12038
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14476 3466 14504 15302
rect 14844 15162 14872 15846
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14568 12918 14596 13670
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14568 11898 14596 12854
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14752 12170 14780 12310
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 11762 14688 12038
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14844 11642 14872 14350
rect 14936 13326 14964 19672
rect 15304 19378 15332 23462
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 17202 15148 17478
rect 15396 17338 15424 25894
rect 15488 24154 15516 37062
rect 15580 35290 15608 39238
rect 15660 38208 15712 38214
rect 15660 38150 15712 38156
rect 15672 37466 15700 38150
rect 15660 37460 15712 37466
rect 15660 37402 15712 37408
rect 15764 37346 15792 40326
rect 15844 38956 15896 38962
rect 15844 38898 15896 38904
rect 15856 38010 15884 38898
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15672 37318 15792 37346
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15672 27402 15700 37318
rect 15844 33040 15896 33046
rect 15844 32982 15896 32988
rect 15856 32434 15884 32982
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15856 31754 15884 32370
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15948 30682 15976 53382
rect 16132 47122 16160 53926
rect 16408 53582 16436 56200
rect 16776 53582 16804 56200
rect 17144 54262 17172 56200
rect 17132 54256 17184 54262
rect 17132 54198 17184 54204
rect 17512 54194 17540 56200
rect 17500 54188 17552 54194
rect 17500 54130 17552 54136
rect 17776 53984 17828 53990
rect 17776 53926 17828 53932
rect 16396 53576 16448 53582
rect 16396 53518 16448 53524
rect 16764 53576 16816 53582
rect 16764 53518 16816 53524
rect 16212 53440 16264 53446
rect 16212 53382 16264 53388
rect 17224 53440 17276 53446
rect 17224 53382 17276 53388
rect 16120 47116 16172 47122
rect 16120 47058 16172 47064
rect 16028 46504 16080 46510
rect 16028 46446 16080 46452
rect 16040 45082 16068 46446
rect 16028 45076 16080 45082
rect 16028 45018 16080 45024
rect 16224 44538 16252 53382
rect 16396 47184 16448 47190
rect 16396 47126 16448 47132
rect 16408 46714 16436 47126
rect 16764 46980 16816 46986
rect 16764 46922 16816 46928
rect 16948 46980 17000 46986
rect 16948 46922 17000 46928
rect 16396 46708 16448 46714
rect 16396 46650 16448 46656
rect 16580 45892 16632 45898
rect 16580 45834 16632 45840
rect 16396 45076 16448 45082
rect 16396 45018 16448 45024
rect 16212 44532 16264 44538
rect 16212 44474 16264 44480
rect 16212 43852 16264 43858
rect 16212 43794 16264 43800
rect 16028 42560 16080 42566
rect 16028 42502 16080 42508
rect 16040 42158 16068 42502
rect 16028 42152 16080 42158
rect 16080 42112 16160 42140
rect 16028 42094 16080 42100
rect 16132 41414 16160 42112
rect 16040 41386 16160 41414
rect 16224 41414 16252 43794
rect 16224 41386 16344 41414
rect 16040 38894 16068 41386
rect 16212 40384 16264 40390
rect 16212 40326 16264 40332
rect 16028 38888 16080 38894
rect 16028 38830 16080 38836
rect 16224 38826 16252 40326
rect 16212 38820 16264 38826
rect 16212 38762 16264 38768
rect 16316 38418 16344 41386
rect 16408 40594 16436 45018
rect 16592 43722 16620 45834
rect 16776 44198 16804 46922
rect 16856 45484 16908 45490
rect 16856 45426 16908 45432
rect 16868 44402 16896 45426
rect 16856 44396 16908 44402
rect 16856 44338 16908 44344
rect 16764 44192 16816 44198
rect 16764 44134 16816 44140
rect 16580 43716 16632 43722
rect 16580 43658 16632 43664
rect 16592 41478 16620 43658
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16580 41472 16632 41478
rect 16580 41414 16632 41420
rect 16396 40588 16448 40594
rect 16396 40530 16448 40536
rect 16488 40588 16540 40594
rect 16488 40530 16540 40536
rect 16396 39636 16448 39642
rect 16396 39578 16448 39584
rect 16408 39506 16436 39578
rect 16396 39500 16448 39506
rect 16396 39442 16448 39448
rect 16500 38842 16528 40530
rect 16684 40526 16712 43046
rect 16764 42628 16816 42634
rect 16764 42570 16816 42576
rect 16672 40520 16724 40526
rect 16672 40462 16724 40468
rect 16580 39908 16632 39914
rect 16580 39850 16632 39856
rect 16592 39030 16620 39850
rect 16580 39024 16632 39030
rect 16580 38966 16632 38972
rect 16408 38814 16528 38842
rect 16304 38412 16356 38418
rect 16304 38354 16356 38360
rect 16120 38208 16172 38214
rect 16212 38208 16264 38214
rect 16120 38150 16172 38156
rect 16210 38176 16212 38185
rect 16264 38176 16266 38185
rect 16132 37874 16160 38150
rect 16210 38111 16266 38120
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16408 37398 16436 38814
rect 16488 38752 16540 38758
rect 16488 38694 16540 38700
rect 16672 38752 16724 38758
rect 16672 38694 16724 38700
rect 16396 37392 16448 37398
rect 16396 37334 16448 37340
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 16028 36916 16080 36922
rect 16028 36858 16080 36864
rect 16040 36106 16068 36858
rect 16224 36718 16252 37266
rect 16212 36712 16264 36718
rect 16210 36680 16212 36689
rect 16264 36680 16266 36689
rect 16120 36644 16172 36650
rect 16210 36615 16266 36624
rect 16120 36586 16172 36592
rect 16028 36100 16080 36106
rect 16028 36042 16080 36048
rect 15764 30654 15976 30682
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15580 25362 15608 27270
rect 15764 27130 15792 30654
rect 15936 30592 15988 30598
rect 15936 30534 15988 30540
rect 15844 29028 15896 29034
rect 15844 28970 15896 28976
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 15752 25696 15804 25702
rect 15752 25638 15804 25644
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15660 25356 15712 25362
rect 15660 25298 15712 25304
rect 15488 24126 15608 24154
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23118 15516 24006
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15580 21865 15608 24126
rect 15672 22778 15700 25298
rect 15764 24274 15792 25638
rect 15752 24268 15804 24274
rect 15752 24210 15804 24216
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15856 21962 15884 28970
rect 15948 27538 15976 30534
rect 16040 29034 16068 36042
rect 16132 32978 16160 36586
rect 16304 36576 16356 36582
rect 16304 36518 16356 36524
rect 16316 36174 16344 36518
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 16304 35692 16356 35698
rect 16304 35634 16356 35640
rect 16316 35442 16344 35634
rect 16408 35630 16436 37334
rect 16396 35624 16448 35630
rect 16396 35566 16448 35572
rect 16316 35414 16436 35442
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 16212 32836 16264 32842
rect 16212 32778 16264 32784
rect 16224 30598 16252 32778
rect 16316 32230 16344 32914
rect 16304 32224 16356 32230
rect 16304 32166 16356 32172
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 16028 29028 16080 29034
rect 16028 28970 16080 28976
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16316 27606 16344 28698
rect 16408 28694 16436 35414
rect 16500 31958 16528 38694
rect 16580 37936 16632 37942
rect 16580 37878 16632 37884
rect 16592 35154 16620 37878
rect 16684 37126 16712 38694
rect 16776 38554 16804 42570
rect 16856 40928 16908 40934
rect 16856 40870 16908 40876
rect 16868 39098 16896 40870
rect 16856 39092 16908 39098
rect 16856 39034 16908 39040
rect 16764 38548 16816 38554
rect 16764 38490 16816 38496
rect 16960 37777 16988 46922
rect 17236 46714 17264 53382
rect 17408 47252 17460 47258
rect 17408 47194 17460 47200
rect 17316 46912 17368 46918
rect 17316 46854 17368 46860
rect 17224 46708 17276 46714
rect 17224 46650 17276 46656
rect 17224 46368 17276 46374
rect 17224 46310 17276 46316
rect 17236 43450 17264 46310
rect 17224 43444 17276 43450
rect 17224 43386 17276 43392
rect 17224 41812 17276 41818
rect 17224 41754 17276 41760
rect 17040 38888 17092 38894
rect 17040 38830 17092 38836
rect 17052 37806 17080 38830
rect 17236 38418 17264 41754
rect 17328 41274 17356 46854
rect 17420 46510 17448 47194
rect 17788 46986 17816 53926
rect 17880 53582 17908 56200
rect 18248 55214 18276 56200
rect 18248 55186 18368 55214
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18340 53582 18368 55186
rect 18616 54194 18644 56200
rect 18604 54188 18656 54194
rect 18604 54130 18656 54136
rect 18512 53984 18564 53990
rect 18512 53926 18564 53932
rect 17868 53576 17920 53582
rect 17868 53518 17920 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 18420 53508 18472 53514
rect 18420 53450 18472 53456
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17776 46980 17828 46986
rect 17776 46922 17828 46928
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 18432 46578 18460 53450
rect 18524 46578 18552 53926
rect 18984 53582 19012 56200
rect 19352 54262 19380 56200
rect 19340 54256 19392 54262
rect 19340 54198 19392 54204
rect 19616 53984 19668 53990
rect 19616 53926 19668 53932
rect 18972 53576 19024 53582
rect 18972 53518 19024 53524
rect 18696 53440 18748 53446
rect 18696 53382 18748 53388
rect 18708 46714 18736 53382
rect 19628 51074 19656 53926
rect 19720 53106 19748 56200
rect 20088 54262 20116 56200
rect 20076 54256 20128 54262
rect 20076 54198 20128 54204
rect 20456 53582 20484 56200
rect 20628 54052 20680 54058
rect 20628 53994 20680 54000
rect 20444 53576 20496 53582
rect 20444 53518 20496 53524
rect 20076 53440 20128 53446
rect 20076 53382 20128 53388
rect 19708 53100 19760 53106
rect 19708 53042 19760 53048
rect 19800 52896 19852 52902
rect 19800 52838 19852 52844
rect 19628 51046 19748 51074
rect 18696 46708 18748 46714
rect 18696 46650 18748 46656
rect 18880 46640 18932 46646
rect 18880 46582 18932 46588
rect 18420 46572 18472 46578
rect 18420 46514 18472 46520
rect 18512 46572 18564 46578
rect 18512 46514 18564 46520
rect 17408 46504 17460 46510
rect 18432 46481 18460 46514
rect 18696 46504 18748 46510
rect 17408 46446 17460 46452
rect 18418 46472 18474 46481
rect 17420 46170 17448 46446
rect 18696 46446 18748 46452
rect 18418 46407 18474 46416
rect 17868 46368 17920 46374
rect 17868 46310 17920 46316
rect 17408 46164 17460 46170
rect 17408 46106 17460 46112
rect 17592 46028 17644 46034
rect 17592 45970 17644 45976
rect 17408 44192 17460 44198
rect 17408 44134 17460 44140
rect 17420 43246 17448 44134
rect 17604 43994 17632 45970
rect 17592 43988 17644 43994
rect 17592 43930 17644 43936
rect 17500 43648 17552 43654
rect 17500 43590 17552 43596
rect 17512 43314 17540 43590
rect 17500 43308 17552 43314
rect 17500 43250 17552 43256
rect 17408 43240 17460 43246
rect 17408 43182 17460 43188
rect 17500 42560 17552 42566
rect 17500 42502 17552 42508
rect 17316 41268 17368 41274
rect 17316 41210 17368 41216
rect 17512 39846 17540 42502
rect 17500 39840 17552 39846
rect 17500 39782 17552 39788
rect 17604 39506 17632 43930
rect 17684 43308 17736 43314
rect 17684 43250 17736 43256
rect 17696 40730 17724 43250
rect 17880 42770 17908 46310
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18512 45552 18564 45558
rect 18512 45494 18564 45500
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 18524 44470 18552 45494
rect 18708 45422 18736 46446
rect 18696 45416 18748 45422
rect 18696 45358 18748 45364
rect 18604 45280 18656 45286
rect 18604 45222 18656 45228
rect 18512 44464 18564 44470
rect 18512 44406 18564 44412
rect 18420 44192 18472 44198
rect 18420 44134 18472 44140
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17868 42764 17920 42770
rect 17868 42706 17920 42712
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 17684 40724 17736 40730
rect 17684 40666 17736 40672
rect 17684 40384 17736 40390
rect 17684 40326 17736 40332
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17408 39432 17460 39438
rect 17408 39374 17460 39380
rect 17316 39024 17368 39030
rect 17316 38966 17368 38972
rect 17224 38412 17276 38418
rect 17224 38354 17276 38360
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 17040 37800 17092 37806
rect 16946 37768 17002 37777
rect 16764 37732 16816 37738
rect 17040 37742 17092 37748
rect 16946 37703 17002 37712
rect 16764 37674 16816 37680
rect 16672 37120 16724 37126
rect 16672 37062 16724 37068
rect 16776 36310 16804 37674
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16856 36848 16908 36854
rect 16856 36790 16908 36796
rect 16764 36304 16816 36310
rect 16764 36246 16816 36252
rect 16868 35834 16896 36790
rect 16856 35828 16908 35834
rect 16856 35770 16908 35776
rect 16580 35148 16632 35154
rect 16580 35090 16632 35096
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16592 32910 16620 33798
rect 16868 32978 16896 34546
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16764 32496 16816 32502
rect 16762 32464 16764 32473
rect 16816 32464 16818 32473
rect 16762 32399 16818 32408
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16488 31952 16540 31958
rect 16488 31894 16540 31900
rect 16776 31686 16804 32302
rect 16868 31890 16896 32914
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 16486 29064 16542 29073
rect 16486 28999 16542 29008
rect 16500 28762 16528 28999
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16396 28688 16448 28694
rect 16396 28630 16448 28636
rect 16304 27600 16356 27606
rect 16304 27542 16356 27548
rect 15936 27532 15988 27538
rect 15936 27474 15988 27480
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 16028 27328 16080 27334
rect 16026 27296 16028 27305
rect 16080 27296 16082 27305
rect 16026 27231 16082 27240
rect 16040 27062 16068 27231
rect 16028 27056 16080 27062
rect 16028 26998 16080 27004
rect 16028 26580 16080 26586
rect 16028 26522 16080 26528
rect 16040 26314 16068 26522
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15936 24812 15988 24818
rect 16040 24800 16068 26250
rect 15988 24772 16068 24800
rect 15936 24754 15988 24760
rect 15948 22710 15976 24754
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15566 21856 15622 21865
rect 15566 21791 15622 21800
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 15632 15068 15638
rect 15016 15574 15068 15580
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14936 11898 14964 12378
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14568 11614 14872 11642
rect 14568 6866 14596 11614
rect 15028 11014 15056 15574
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14752 3398 14780 10950
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14844 3058 14872 9862
rect 15120 6914 15148 17138
rect 15488 16658 15516 17682
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15382 16552 15438 16561
rect 15382 16487 15438 16496
rect 15198 16280 15254 16289
rect 15198 16215 15254 16224
rect 15212 12170 15240 16215
rect 15396 16114 15424 16487
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15488 16046 15516 16594
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15304 15094 15332 15982
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15304 12986 15332 14282
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15488 11694 15516 15982
rect 15580 14006 15608 21791
rect 15856 21622 15884 21898
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19394 15884 20198
rect 15948 19514 15976 22374
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16040 20806 16068 21898
rect 16132 21894 16160 27338
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16224 24750 16252 26522
rect 16408 26330 16436 28630
rect 16580 27872 16632 27878
rect 16580 27814 16632 27820
rect 16408 26302 16528 26330
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16408 25838 16436 26182
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16316 24750 16344 25162
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16224 24274 16252 24686
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16118 21720 16174 21729
rect 16118 21655 16174 21664
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 20398 16068 20742
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15856 19366 15976 19394
rect 15948 18630 15976 19366
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 14226 15700 16390
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15672 14198 15792 14226
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15672 12850 15700 13942
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 11830 15700 12786
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 15028 6886 15148 6914
rect 15028 3126 15056 6886
rect 15212 4146 15240 9386
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14384 800 14412 2450
rect 14752 800 14780 2926
rect 15304 2650 15332 11630
rect 15764 11150 15792 14198
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 8634 15792 11086
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15856 5642 15884 15030
rect 15948 8974 15976 18566
rect 16132 16182 16160 21655
rect 16224 16590 16252 23190
rect 16316 23186 16344 24686
rect 16408 23662 16436 25774
rect 16500 23730 16528 26302
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16304 23180 16356 23186
rect 16304 23122 16356 23128
rect 16408 22778 16436 23598
rect 16592 23118 16620 27814
rect 16684 25158 16712 30534
rect 16868 30410 16896 31826
rect 16776 30382 16896 30410
rect 16960 30394 16988 37062
rect 17052 35766 17080 37742
rect 17144 36786 17172 38150
rect 17236 37398 17264 38354
rect 17224 37392 17276 37398
rect 17224 37334 17276 37340
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17040 35760 17092 35766
rect 17328 35714 17356 38966
rect 17040 35702 17092 35708
rect 17052 34678 17080 35702
rect 17236 35686 17356 35714
rect 17132 35556 17184 35562
rect 17132 35498 17184 35504
rect 17144 35222 17172 35498
rect 17132 35216 17184 35222
rect 17132 35158 17184 35164
rect 17040 34672 17092 34678
rect 17040 34614 17092 34620
rect 17132 34536 17184 34542
rect 17132 34478 17184 34484
rect 17144 34202 17172 34478
rect 17132 34196 17184 34202
rect 17132 34138 17184 34144
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 17052 32774 17080 33934
rect 17132 33584 17184 33590
rect 17132 33526 17184 33532
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17052 32298 17080 32710
rect 17040 32292 17092 32298
rect 17040 32234 17092 32240
rect 17038 32192 17094 32201
rect 17038 32127 17094 32136
rect 17052 30954 17080 32127
rect 17144 31482 17172 33526
rect 17236 32042 17264 35686
rect 17316 35624 17368 35630
rect 17316 35566 17368 35572
rect 17328 35290 17356 35566
rect 17316 35284 17368 35290
rect 17316 35226 17368 35232
rect 17314 32600 17370 32609
rect 17314 32535 17316 32544
rect 17368 32535 17370 32544
rect 17316 32506 17368 32512
rect 17420 32502 17448 39374
rect 17592 39364 17644 39370
rect 17592 39306 17644 39312
rect 17604 38282 17632 39306
rect 17592 38276 17644 38282
rect 17592 38218 17644 38224
rect 17592 37120 17644 37126
rect 17590 37088 17592 37097
rect 17644 37088 17646 37097
rect 17590 37023 17646 37032
rect 17696 36854 17724 40326
rect 17788 39352 17816 42502
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17868 42220 17920 42226
rect 17868 42162 17920 42168
rect 17880 41682 17908 42162
rect 17868 41676 17920 41682
rect 17868 41618 17920 41624
rect 18328 41472 18380 41478
rect 18328 41414 18380 41420
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 17880 39982 17908 40666
rect 18340 40526 18368 41414
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18328 40384 18380 40390
rect 18432 40372 18460 44134
rect 18524 42276 18552 44406
rect 18616 43858 18644 45222
rect 18708 44538 18736 45358
rect 18696 44532 18748 44538
rect 18696 44474 18748 44480
rect 18604 43852 18656 43858
rect 18604 43794 18656 43800
rect 18616 42838 18644 43794
rect 18788 43784 18840 43790
rect 18788 43726 18840 43732
rect 18604 42832 18656 42838
rect 18604 42774 18656 42780
rect 18604 42288 18656 42294
rect 18524 42248 18604 42276
rect 18524 41546 18552 42248
rect 18604 42230 18656 42236
rect 18604 42152 18656 42158
rect 18604 42094 18656 42100
rect 18512 41540 18564 41546
rect 18512 41482 18564 41488
rect 18524 40934 18552 41482
rect 18512 40928 18564 40934
rect 18512 40870 18564 40876
rect 18616 40594 18644 42094
rect 18800 41682 18828 43726
rect 18788 41676 18840 41682
rect 18788 41618 18840 41624
rect 18800 41206 18828 41618
rect 18788 41200 18840 41206
rect 18788 41142 18840 41148
rect 18696 41064 18748 41070
rect 18696 41006 18748 41012
rect 18604 40588 18656 40594
rect 18604 40530 18656 40536
rect 18512 40520 18564 40526
rect 18512 40462 18564 40468
rect 18380 40344 18460 40372
rect 18328 40326 18380 40332
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17868 39976 17920 39982
rect 17868 39918 17920 39924
rect 18052 39840 18104 39846
rect 18052 39782 18104 39788
rect 18064 39506 18092 39782
rect 18052 39500 18104 39506
rect 18052 39442 18104 39448
rect 17960 39364 18012 39370
rect 17788 39324 17960 39352
rect 17684 36848 17736 36854
rect 17684 36790 17736 36796
rect 17500 36780 17552 36786
rect 17500 36722 17552 36728
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 17408 32292 17460 32298
rect 17408 32234 17460 32240
rect 17236 32014 17356 32042
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 17052 30926 17172 30954
rect 17040 30864 17092 30870
rect 17040 30806 17092 30812
rect 16948 30388 17000 30394
rect 16776 29034 16804 30382
rect 16948 30330 17000 30336
rect 16948 30184 17000 30190
rect 16948 30126 17000 30132
rect 16960 29050 16988 30126
rect 16764 29028 16816 29034
rect 16764 28970 16816 28976
rect 16868 29022 16988 29050
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16776 26586 16804 27950
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 16868 26314 16896 29022
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16960 27470 16988 28358
rect 17052 27538 17080 30806
rect 17144 29238 17172 30926
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17040 27532 17092 27538
rect 17040 27474 17092 27480
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 17144 27282 17172 29174
rect 17236 27538 17264 31894
rect 17328 30802 17356 32014
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17420 30734 17448 32234
rect 17512 31958 17540 36722
rect 17590 36544 17646 36553
rect 17590 36479 17646 36488
rect 17604 36106 17632 36479
rect 17682 36408 17738 36417
rect 17682 36343 17738 36352
rect 17696 36242 17724 36343
rect 17684 36236 17736 36242
rect 17684 36178 17736 36184
rect 17788 36122 17816 39324
rect 17960 39306 18012 39312
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17868 37800 17920 37806
rect 17866 37768 17868 37777
rect 17920 37768 17922 37777
rect 17866 37703 17922 37712
rect 18052 37664 18104 37670
rect 18052 37606 18104 37612
rect 18064 37330 18092 37606
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 18340 36922 18368 40326
rect 18420 39840 18472 39846
rect 18420 39782 18472 39788
rect 18432 39030 18460 39782
rect 18420 39024 18472 39030
rect 18420 38966 18472 38972
rect 18432 37874 18460 38966
rect 18420 37868 18472 37874
rect 18420 37810 18472 37816
rect 18524 37670 18552 40462
rect 18604 40452 18656 40458
rect 18604 40394 18656 40400
rect 18616 39098 18644 40394
rect 18604 39092 18656 39098
rect 18604 39034 18656 39040
rect 18604 38276 18656 38282
rect 18604 38218 18656 38224
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18512 36712 18564 36718
rect 18326 36680 18382 36689
rect 18510 36680 18512 36689
rect 18564 36680 18566 36689
rect 18326 36615 18382 36624
rect 18420 36644 18472 36650
rect 17592 36100 17644 36106
rect 17592 36042 17644 36048
rect 17696 36094 17816 36122
rect 17592 32292 17644 32298
rect 17592 32234 17644 32240
rect 17500 31952 17552 31958
rect 17500 31894 17552 31900
rect 17408 30728 17460 30734
rect 17408 30670 17460 30676
rect 17604 30190 17632 32234
rect 17696 32201 17724 36094
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17960 35216 18012 35222
rect 17960 35158 18012 35164
rect 17972 34932 18000 35158
rect 17880 34904 18000 34932
rect 17880 34728 17908 34904
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17880 34700 18000 34728
rect 17972 33998 18000 34700
rect 18340 34542 18368 36615
rect 18510 36615 18566 36624
rect 18420 36586 18472 36592
rect 18328 34536 18380 34542
rect 18328 34478 18380 34484
rect 18432 34066 18460 36586
rect 18616 36378 18644 38218
rect 18604 36372 18656 36378
rect 18604 36314 18656 36320
rect 18708 36310 18736 41006
rect 18788 40928 18840 40934
rect 18788 40870 18840 40876
rect 18800 39846 18828 40870
rect 18788 39840 18840 39846
rect 18788 39782 18840 39788
rect 18788 39636 18840 39642
rect 18788 39578 18840 39584
rect 18800 38010 18828 39578
rect 18788 38004 18840 38010
rect 18788 37946 18840 37952
rect 18696 36304 18748 36310
rect 18696 36246 18748 36252
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18432 32434 18460 34002
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 17776 32224 17828 32230
rect 17682 32192 17738 32201
rect 17776 32166 17828 32172
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 17682 32127 17738 32136
rect 17788 31890 17816 32166
rect 17776 31884 17828 31890
rect 17776 31826 17828 31832
rect 17868 31884 17920 31890
rect 17868 31826 17920 31832
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 17592 30184 17644 30190
rect 17592 30126 17644 30132
rect 17316 30048 17368 30054
rect 17316 29990 17368 29996
rect 17328 28218 17356 29990
rect 17500 29504 17552 29510
rect 17592 29504 17644 29510
rect 17500 29446 17552 29452
rect 17590 29472 17592 29481
rect 17644 29472 17646 29481
rect 17512 29306 17540 29446
rect 17590 29407 17646 29416
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17420 28218 17448 28358
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 16960 27254 17172 27282
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 25974 16804 26182
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16670 24848 16726 24857
rect 16670 24783 16726 24792
rect 16684 24206 16712 24783
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16500 21962 16528 22646
rect 16684 22094 16712 24142
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16776 22574 16804 22918
rect 16868 22642 16896 25230
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16684 22066 16804 22094
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16500 20874 16528 21898
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 18766 16620 20742
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 18086 16620 18566
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 14006 16068 14282
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16040 11082 16068 13398
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 16040 8786 16068 11018
rect 15948 8758 16068 8786
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15120 800 15148 2450
rect 15488 800 15516 3538
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15856 800 15884 2926
rect 15948 2582 15976 8758
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16040 6798 16068 8570
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 3670 16068 5170
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16132 3534 16160 13194
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16224 11626 16252 12786
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16224 800 16252 4014
rect 16316 2446 16344 15914
rect 16592 12442 16620 18022
rect 16684 17882 16712 21082
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16776 15502 16804 22066
rect 16868 22080 16896 22578
rect 16960 22273 16988 27254
rect 17236 27010 17264 27270
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17052 26982 17264 27010
rect 16946 22264 17002 22273
rect 16946 22199 17002 22208
rect 16948 22092 17000 22098
rect 16868 22052 16948 22080
rect 16948 22034 17000 22040
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16960 20602 16988 20878
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17052 20466 17080 26982
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17144 22438 17172 26794
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17316 26240 17368 26246
rect 17316 26182 17368 26188
rect 17328 24596 17356 26182
rect 17420 24750 17448 26726
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17328 24568 17448 24596
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 17130 22264 17186 22273
rect 17130 22199 17186 22208
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17040 19440 17092 19446
rect 17038 19408 17040 19417
rect 17092 19408 17094 19417
rect 17038 19343 17094 19352
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16868 14482 16896 16050
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 13938 16896 14418
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16408 11150 16436 12310
rect 16500 11370 16528 12378
rect 16500 11342 16620 11370
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16592 7886 16620 11342
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16684 3058 16712 13806
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16592 800 16620 2858
rect 16776 2446 16804 12106
rect 16868 11762 16896 13874
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16960 800 16988 2382
rect 17052 2378 17080 19110
rect 17144 18834 17172 22199
rect 17236 22030 17264 22918
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17328 21554 17356 22918
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17314 20632 17370 20641
rect 17420 20602 17448 24568
rect 17512 22137 17540 27066
rect 17696 24274 17724 31282
rect 17880 29050 17908 31826
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18144 29096 18196 29102
rect 17880 29044 18144 29050
rect 17880 29038 18196 29044
rect 17880 29022 18184 29038
rect 17880 28626 17908 29022
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18340 28200 18368 29514
rect 18248 28172 18368 28200
rect 17958 27568 18014 27577
rect 17958 27503 18014 27512
rect 17972 27470 18000 27503
rect 17960 27464 18012 27470
rect 17866 27432 17922 27441
rect 17960 27406 18012 27412
rect 18248 27418 18276 28172
rect 18432 28098 18460 32166
rect 18524 30326 18552 35974
rect 18604 35828 18656 35834
rect 18604 35770 18656 35776
rect 18616 35737 18644 35770
rect 18800 35766 18828 37946
rect 18892 36689 18920 46582
rect 19616 45824 19668 45830
rect 19720 45812 19748 51046
rect 19812 46034 19840 52838
rect 19800 46028 19852 46034
rect 19800 45970 19852 45976
rect 19984 46028 20036 46034
rect 19984 45970 20036 45976
rect 19800 45824 19852 45830
rect 19720 45792 19800 45812
rect 19852 45792 19854 45801
rect 19720 45784 19798 45792
rect 19616 45766 19668 45772
rect 19156 45552 19208 45558
rect 19156 45494 19208 45500
rect 19064 41744 19116 41750
rect 19064 41686 19116 41692
rect 19076 41070 19104 41686
rect 19064 41064 19116 41070
rect 19064 41006 19116 41012
rect 19064 40656 19116 40662
rect 19064 40598 19116 40604
rect 18972 39296 19024 39302
rect 18972 39238 19024 39244
rect 18878 36680 18934 36689
rect 18878 36615 18934 36624
rect 18788 35760 18840 35766
rect 18602 35728 18658 35737
rect 18788 35702 18840 35708
rect 18602 35663 18658 35672
rect 18984 35222 19012 39238
rect 19076 39080 19104 40598
rect 19168 40089 19196 45494
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 19340 44736 19392 44742
rect 19340 44678 19392 44684
rect 19352 42158 19380 44678
rect 19444 42770 19472 44814
rect 19524 44328 19576 44334
rect 19524 44270 19576 44276
rect 19432 42764 19484 42770
rect 19432 42706 19484 42712
rect 19536 42362 19564 44270
rect 19524 42356 19576 42362
rect 19524 42298 19576 42304
rect 19432 42220 19484 42226
rect 19432 42162 19484 42168
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 19444 41614 19472 42162
rect 19432 41608 19484 41614
rect 19432 41550 19484 41556
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 19248 41200 19300 41206
rect 19248 41142 19300 41148
rect 19260 40934 19288 41142
rect 19248 40928 19300 40934
rect 19248 40870 19300 40876
rect 19154 40080 19210 40089
rect 19154 40015 19210 40024
rect 19248 39568 19300 39574
rect 19248 39510 19300 39516
rect 19076 39052 19196 39080
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19076 36106 19104 37810
rect 19064 36100 19116 36106
rect 19064 36042 19116 36048
rect 18972 35216 19024 35222
rect 18972 35158 19024 35164
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18708 31754 18736 34954
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 18696 31748 18748 31754
rect 18696 31690 18748 31696
rect 18788 31204 18840 31210
rect 18788 31146 18840 31152
rect 18512 30320 18564 30326
rect 18512 30262 18564 30268
rect 18604 30320 18656 30326
rect 18604 30262 18656 30268
rect 18512 30116 18564 30122
rect 18512 30058 18564 30064
rect 18340 28082 18460 28098
rect 18328 28076 18460 28082
rect 18380 28070 18460 28076
rect 18328 28018 18380 28024
rect 18420 28008 18472 28014
rect 18418 27976 18420 27985
rect 18472 27976 18474 27985
rect 18418 27911 18474 27920
rect 18418 27568 18474 27577
rect 18524 27538 18552 30058
rect 18616 28966 18644 30262
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 28014 18644 28902
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18418 27503 18420 27512
rect 18472 27503 18474 27512
rect 18512 27532 18564 27538
rect 18420 27474 18472 27480
rect 18512 27474 18564 27480
rect 18248 27390 18368 27418
rect 17866 27367 17922 27376
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17788 26450 17816 27270
rect 17880 27130 17908 27367
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17868 27124 17920 27130
rect 17868 27066 17920 27072
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17788 25838 17816 26386
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17880 24070 17908 25910
rect 18340 25362 18368 27390
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17590 23488 17646 23497
rect 17590 23423 17646 23432
rect 17604 22574 17632 23423
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17498 22128 17554 22137
rect 17498 22063 17554 22072
rect 17512 21690 17540 22063
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17314 20567 17370 20576
rect 17408 20596 17460 20602
rect 17222 20496 17278 20505
rect 17222 20431 17278 20440
rect 17236 19446 17264 20431
rect 17328 19854 17356 20567
rect 17408 20538 17460 20544
rect 17512 20482 17540 20810
rect 17420 20454 17540 20482
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17420 19700 17448 20454
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17328 19672 17448 19700
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17328 17678 17356 19672
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17420 17746 17448 18158
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 17270 17356 17614
rect 17316 17264 17368 17270
rect 17316 17206 17368 17212
rect 17420 17202 17448 17682
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17144 16046 17172 17070
rect 17420 16182 17448 17138
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 14618 17172 15982
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17132 13864 17184 13870
rect 17236 13852 17264 14826
rect 17420 14362 17448 15370
rect 17512 14940 17540 19722
rect 17604 18170 17632 22510
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17696 22166 17724 22374
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17788 22098 17816 24006
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17880 22001 17908 24006
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17866 21992 17922 22001
rect 17866 21927 17922 21936
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17880 20942 17908 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 19718 18276 20198
rect 18340 19854 18368 21558
rect 18432 19922 18460 24550
rect 18524 24274 18552 27474
rect 18616 27402 18644 27950
rect 18604 27396 18656 27402
rect 18604 27338 18656 27344
rect 18708 26926 18736 29582
rect 18800 27062 18828 31146
rect 18892 29050 18920 34886
rect 19076 34678 19104 36042
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 18972 33924 19024 33930
rect 18972 33866 19024 33872
rect 18984 33522 19012 33866
rect 18972 33516 19024 33522
rect 18972 33458 19024 33464
rect 18972 33040 19024 33046
rect 18972 32982 19024 32988
rect 18984 32366 19012 32982
rect 19076 32842 19104 34614
rect 19168 32910 19196 39052
rect 19260 36922 19288 39510
rect 19352 38418 19380 41414
rect 19340 38412 19392 38418
rect 19340 38354 19392 38360
rect 19444 37942 19472 41550
rect 19524 41472 19576 41478
rect 19524 41414 19576 41420
rect 19536 39642 19564 41414
rect 19628 40594 19656 45766
rect 19798 45727 19854 45736
rect 19708 45280 19760 45286
rect 19708 45222 19760 45228
rect 19720 41682 19748 45222
rect 19996 44810 20024 45970
rect 20088 45558 20116 53382
rect 20640 45830 20668 53994
rect 20824 53582 20852 56200
rect 21192 54194 21220 56200
rect 21180 54188 21232 54194
rect 21180 54130 21232 54136
rect 20996 53984 21048 53990
rect 20996 53926 21048 53932
rect 20812 53576 20864 53582
rect 20812 53518 20864 53524
rect 21008 51074 21036 53926
rect 21560 53582 21588 56200
rect 21824 53984 21876 53990
rect 21824 53926 21876 53932
rect 21548 53576 21600 53582
rect 21548 53518 21600 53524
rect 21456 53440 21508 53446
rect 21456 53382 21508 53388
rect 21548 53440 21600 53446
rect 21548 53382 21600 53388
rect 21468 51074 21496 53382
rect 21008 51046 21128 51074
rect 20628 45824 20680 45830
rect 20628 45766 20680 45772
rect 20640 45665 20668 45766
rect 20626 45656 20682 45665
rect 20626 45591 20682 45600
rect 20076 45552 20128 45558
rect 20076 45494 20128 45500
rect 20352 45416 20404 45422
rect 20352 45358 20404 45364
rect 19800 44804 19852 44810
rect 19800 44746 19852 44752
rect 19984 44804 20036 44810
rect 19984 44746 20036 44752
rect 19812 43994 19840 44746
rect 20364 44198 20392 45358
rect 20996 44804 21048 44810
rect 20996 44746 21048 44752
rect 20904 44532 20956 44538
rect 20904 44474 20956 44480
rect 20352 44192 20404 44198
rect 20352 44134 20404 44140
rect 19800 43988 19852 43994
rect 19800 43930 19852 43936
rect 20076 43852 20128 43858
rect 20076 43794 20128 43800
rect 19708 41676 19760 41682
rect 19708 41618 19760 41624
rect 20088 40934 20116 43794
rect 20364 42906 20392 44134
rect 20352 42900 20404 42906
rect 20352 42842 20404 42848
rect 20260 41744 20312 41750
rect 20260 41686 20312 41692
rect 20076 40928 20128 40934
rect 20076 40870 20128 40876
rect 19616 40588 19668 40594
rect 19616 40530 19668 40536
rect 19708 40384 19760 40390
rect 19708 40326 19760 40332
rect 19616 39976 19668 39982
rect 19616 39918 19668 39924
rect 19524 39636 19576 39642
rect 19524 39578 19576 39584
rect 19628 39370 19656 39918
rect 19616 39364 19668 39370
rect 19616 39306 19668 39312
rect 19720 39098 19748 40326
rect 19892 39296 19944 39302
rect 19944 39256 20024 39284
rect 19892 39238 19944 39244
rect 19708 39092 19760 39098
rect 19708 39034 19760 39040
rect 19616 38820 19668 38826
rect 19616 38762 19668 38768
rect 19524 38752 19576 38758
rect 19524 38694 19576 38700
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 19340 37392 19392 37398
rect 19340 37334 19392 37340
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19248 36100 19300 36106
rect 19248 36042 19300 36048
rect 19260 35748 19288 36042
rect 19352 36038 19380 37334
rect 19444 37194 19472 37878
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19444 36786 19472 37130
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19340 35760 19392 35766
rect 19260 35720 19340 35748
rect 19340 35702 19392 35708
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 19260 34542 19288 35566
rect 19340 35488 19392 35494
rect 19340 35430 19392 35436
rect 19352 35222 19380 35430
rect 19536 35306 19564 38694
rect 19628 38010 19656 38762
rect 19996 38282 20024 39256
rect 20088 38418 20116 40870
rect 20272 40118 20300 41686
rect 20260 40112 20312 40118
rect 20260 40054 20312 40060
rect 20076 38412 20128 38418
rect 20076 38354 20128 38360
rect 20272 38298 20300 40054
rect 20364 39506 20392 42842
rect 20444 42356 20496 42362
rect 20444 42298 20496 42304
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20456 38894 20484 42298
rect 20720 42220 20772 42226
rect 20720 42162 20772 42168
rect 20536 39908 20588 39914
rect 20536 39850 20588 39856
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 19984 38276 20036 38282
rect 19984 38218 20036 38224
rect 20088 38270 20300 38298
rect 19616 38004 19668 38010
rect 19668 37964 19748 37992
rect 19616 37946 19668 37952
rect 19616 37664 19668 37670
rect 19616 37606 19668 37612
rect 19628 37262 19656 37606
rect 19616 37256 19668 37262
rect 19616 37198 19668 37204
rect 19720 36718 19748 37964
rect 19800 36848 19852 36854
rect 19800 36790 19852 36796
rect 19708 36712 19760 36718
rect 19708 36654 19760 36660
rect 19444 35278 19564 35306
rect 19708 35284 19760 35290
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19248 34536 19300 34542
rect 19248 34478 19300 34484
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 19064 32836 19116 32842
rect 19064 32778 19116 32784
rect 18972 32360 19024 32366
rect 18972 32302 19024 32308
rect 18984 30326 19012 32302
rect 18972 30320 19024 30326
rect 18972 30262 19024 30268
rect 18972 29504 19024 29510
rect 18972 29446 19024 29452
rect 18984 29345 19012 29446
rect 18970 29336 19026 29345
rect 18970 29271 19026 29280
rect 19076 29238 19104 32778
rect 19352 32570 19380 35158
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19154 30288 19210 30297
rect 19154 30223 19156 30232
rect 19208 30223 19210 30232
rect 19156 30194 19208 30200
rect 19064 29232 19116 29238
rect 19064 29174 19116 29180
rect 18892 29034 19104 29050
rect 18892 29028 19116 29034
rect 18892 29022 19064 29028
rect 18892 28150 18920 29022
rect 19064 28970 19116 28976
rect 18880 28144 18932 28150
rect 18880 28086 18932 28092
rect 18878 27976 18934 27985
rect 18878 27911 18934 27920
rect 18788 27056 18840 27062
rect 18788 26998 18840 27004
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18524 23186 18552 24210
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18616 22794 18644 24686
rect 18524 22778 18644 22794
rect 18512 22772 18644 22778
rect 18564 22766 18644 22772
rect 18512 22714 18564 22720
rect 18524 20398 18552 22714
rect 18708 22556 18736 25638
rect 18892 24138 18920 27911
rect 19064 25220 19116 25226
rect 19064 25162 19116 25168
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18616 22528 18736 22556
rect 18616 21010 18644 22528
rect 18800 22094 18828 24006
rect 18892 23322 18920 24074
rect 18880 23316 18932 23322
rect 18880 23258 18932 23264
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 22438 18920 23122
rect 19076 22710 19104 25162
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18984 22234 19012 22510
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19076 22234 19104 22374
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18708 22066 18828 22094
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18340 18358 18368 19790
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 17604 18142 17908 18170
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 15502 17816 16934
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17880 15042 17908 18142
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18156 16454 18184 17206
rect 18340 16590 18368 18294
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18432 17338 18460 17750
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18340 16046 18368 16390
rect 18432 16250 18460 17070
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15450 18368 15982
rect 18432 15570 18460 16186
rect 18524 15638 18552 18702
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18340 15422 18460 15450
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17880 15014 18000 15042
rect 17512 14912 17908 14940
rect 17420 14334 17540 14362
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17184 13824 17264 13852
rect 17132 13806 17184 13812
rect 17144 11898 17172 13806
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17236 12986 17264 13262
rect 17328 12986 17356 14010
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17420 11830 17448 14214
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17420 6914 17448 11766
rect 17328 6886 17448 6914
rect 17328 6322 17356 6886
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17512 4622 17540 14334
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 17328 800 17356 2790
rect 17696 800 17724 3538
rect 17788 3534 17816 8842
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17880 3058 17908 14912
rect 17972 14346 18000 15014
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 13394 18368 14758
rect 18432 14074 18460 15422
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18524 15026 18552 15302
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18616 14414 18644 19722
rect 18708 19378 18736 22066
rect 18984 21622 19012 22170
rect 18972 21616 19024 21622
rect 18972 21558 19024 21564
rect 18984 21010 19012 21558
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18984 20534 19012 20946
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18786 19408 18842 19417
rect 18696 19372 18748 19378
rect 18786 19343 18842 19352
rect 18696 19314 18748 19320
rect 18800 17882 18828 19343
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18290 19012 19110
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18708 14074 18736 17546
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10742 18368 12854
rect 18432 12102 18460 13874
rect 18708 13394 18736 14010
rect 18800 13938 18828 17682
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18800 13326 18828 13670
rect 18892 13462 18920 15302
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12986 18552 13126
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18984 12434 19012 18226
rect 19076 15162 19104 18634
rect 19168 17678 19196 30194
rect 19248 29844 19300 29850
rect 19248 29786 19300 29792
rect 19260 28014 19288 29786
rect 19352 29714 19380 32166
rect 19444 31414 19472 35278
rect 19708 35226 19760 35232
rect 19616 35148 19668 35154
rect 19616 35090 19668 35096
rect 19522 34640 19578 34649
rect 19522 34575 19578 34584
rect 19536 34542 19564 34575
rect 19524 34536 19576 34542
rect 19524 34478 19576 34484
rect 19628 33046 19656 35090
rect 19616 33040 19668 33046
rect 19616 32982 19668 32988
rect 19720 32570 19748 35226
rect 19812 33862 19840 36790
rect 19996 35170 20024 38218
rect 19904 35142 20024 35170
rect 19904 34134 19932 35142
rect 20088 35018 20116 38270
rect 20260 38208 20312 38214
rect 20260 38150 20312 38156
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 20180 35834 20208 37130
rect 20168 35828 20220 35834
rect 20168 35770 20220 35776
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 19892 34128 19944 34134
rect 19892 34070 19944 34076
rect 19800 33856 19852 33862
rect 19800 33798 19852 33804
rect 19984 33448 20036 33454
rect 20036 33408 20116 33436
rect 19984 33390 20036 33396
rect 19708 32564 19760 32570
rect 19708 32506 19760 32512
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 19708 31680 19760 31686
rect 19708 31622 19760 31628
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 19432 30116 19484 30122
rect 19432 30058 19484 30064
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19352 24954 19380 29446
rect 19444 28082 19472 30058
rect 19616 29776 19668 29782
rect 19616 29718 19668 29724
rect 19522 29336 19578 29345
rect 19522 29271 19524 29280
rect 19576 29271 19578 29280
rect 19524 29242 19576 29248
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 19536 26042 19564 27542
rect 19628 27062 19656 29718
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19444 24818 19472 25978
rect 19628 25838 19656 26998
rect 19720 26926 19748 31622
rect 19892 30320 19944 30326
rect 19892 30262 19944 30268
rect 19904 29492 19932 30262
rect 19996 29510 20024 31962
rect 20088 31686 20116 33408
rect 20168 33380 20220 33386
rect 20168 33322 20220 33328
rect 20180 31754 20208 33322
rect 20272 32434 20300 38150
rect 20548 37890 20576 39850
rect 20732 39642 20760 42162
rect 20812 41268 20864 41274
rect 20812 41210 20864 41216
rect 20720 39636 20772 39642
rect 20720 39578 20772 39584
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20640 38196 20668 39238
rect 20720 38208 20772 38214
rect 20640 38168 20720 38196
rect 20720 38150 20772 38156
rect 20456 37862 20576 37890
rect 20456 36281 20484 37862
rect 20536 37732 20588 37738
rect 20536 37674 20588 37680
rect 20442 36272 20498 36281
rect 20442 36207 20498 36216
rect 20350 36136 20406 36145
rect 20350 36071 20352 36080
rect 20404 36071 20406 36080
rect 20352 36042 20404 36048
rect 20548 34066 20576 37674
rect 20732 37369 20760 38150
rect 20718 37360 20774 37369
rect 20718 37295 20774 37304
rect 20720 36644 20772 36650
rect 20720 36586 20772 36592
rect 20628 36576 20680 36582
rect 20732 36553 20760 36586
rect 20628 36518 20680 36524
rect 20718 36544 20774 36553
rect 20640 36242 20668 36518
rect 20718 36479 20774 36488
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20626 36136 20682 36145
rect 20626 36071 20682 36080
rect 20536 34060 20588 34066
rect 20456 34020 20536 34048
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20364 33454 20392 33934
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 20364 32978 20392 33390
rect 20456 33114 20484 34020
rect 20536 34002 20588 34008
rect 20444 33108 20496 33114
rect 20444 33050 20496 33056
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 20350 32736 20406 32745
rect 20350 32671 20406 32680
rect 20260 32428 20312 32434
rect 20260 32370 20312 32376
rect 20364 32026 20392 32671
rect 20640 32314 20668 36071
rect 20824 36038 20852 41210
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20732 35154 20760 35974
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 20732 33658 20760 34954
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20824 33658 20852 33798
rect 20720 33652 20772 33658
rect 20720 33594 20772 33600
rect 20812 33652 20864 33658
rect 20812 33594 20864 33600
rect 20720 32836 20772 32842
rect 20720 32778 20772 32784
rect 20456 32286 20668 32314
rect 20456 32230 20484 32286
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 20536 32224 20588 32230
rect 20536 32166 20588 32172
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20444 31952 20496 31958
rect 20444 31894 20496 31900
rect 20180 31726 20392 31754
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 20166 30288 20222 30297
rect 20166 30223 20168 30232
rect 20220 30223 20222 30232
rect 20168 30194 20220 30200
rect 19812 29464 19932 29492
rect 19984 29504 20036 29510
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19708 25832 19760 25838
rect 19708 25774 19760 25780
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19536 24954 19564 25638
rect 19628 25498 19656 25774
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 19786 19288 22918
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19352 21690 19380 22510
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19352 21078 19380 21626
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19444 20942 19472 24346
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19536 21418 19564 23258
rect 19720 22166 19748 25774
rect 19812 25498 19840 29464
rect 19984 29446 20036 29452
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19892 27872 19944 27878
rect 19892 27814 19944 27820
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19812 24206 19840 24550
rect 19904 24274 19932 27814
rect 19996 26314 20024 28494
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 20088 26926 20116 27950
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19800 24200 19852 24206
rect 19800 24142 19852 24148
rect 19800 22704 19852 22710
rect 19800 22646 19852 22652
rect 19812 22438 19840 22646
rect 20180 22522 20208 30194
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20272 26790 20300 30126
rect 20364 28558 20392 31726
rect 20456 30326 20484 31894
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 20260 26784 20312 26790
rect 20260 26726 20312 26732
rect 20272 26450 20300 26726
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20364 25362 20392 27066
rect 20456 25906 20484 29990
rect 20548 28150 20576 32166
rect 20732 32065 20760 32778
rect 20812 32496 20864 32502
rect 20810 32464 20812 32473
rect 20864 32464 20866 32473
rect 20810 32399 20866 32408
rect 20812 32360 20864 32366
rect 20812 32302 20864 32308
rect 20718 32056 20774 32065
rect 20718 31991 20774 32000
rect 20628 31748 20680 31754
rect 20628 31690 20680 31696
rect 20640 29238 20668 31690
rect 20824 31464 20852 32302
rect 20732 31436 20852 31464
rect 20732 29782 20760 31436
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20824 30326 20852 31282
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20720 29776 20772 29782
rect 20720 29718 20772 29724
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20640 25362 20668 26862
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20640 24750 20668 25298
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20180 22494 20484 22522
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 19708 22160 19760 22166
rect 20076 22160 20128 22166
rect 19708 22102 19760 22108
rect 19798 22128 19854 22137
rect 19616 22092 19668 22098
rect 20128 22108 20208 22114
rect 20076 22102 20208 22108
rect 20088 22086 20208 22102
rect 19798 22063 19854 22072
rect 19616 22034 19668 22040
rect 19628 21554 19656 22034
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19524 21412 19576 21418
rect 19524 21354 19576 21360
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19536 18986 19564 21354
rect 19536 18958 19656 18986
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19260 17746 19288 18770
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19260 17338 19288 17682
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19260 12782 19288 13262
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 18800 12406 19012 12434
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18064 4690 18092 5170
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 18340 2854 18368 4490
rect 18708 4146 18736 12106
rect 18800 8974 18828 12406
rect 19260 10810 19288 12718
rect 19352 12434 19380 17818
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 17338 19472 17614
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15162 19564 15846
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19628 13258 19656 18958
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 13852 19748 17478
rect 19812 14006 19840 22063
rect 20180 21894 20208 22086
rect 20364 21962 20392 22374
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 19904 21622 19932 21830
rect 20364 21622 20392 21898
rect 19892 21616 19944 21622
rect 19892 21558 19944 21564
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20364 20806 20392 21558
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20534 20392 20742
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19890 18864 19946 18873
rect 19890 18799 19892 18808
rect 19944 18799 19946 18808
rect 19892 18770 19944 18776
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19996 17270 20024 17478
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19890 15600 19946 15609
rect 19890 15535 19892 15544
rect 19944 15535 19946 15544
rect 19892 15506 19944 15512
rect 20088 15314 20116 18022
rect 20180 15434 20208 18566
rect 20272 17882 20300 19110
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20364 17746 20392 20470
rect 20456 19174 20484 22494
rect 20640 21570 20668 24006
rect 20732 23322 20760 28562
rect 20824 28422 20852 28698
rect 20916 28626 20944 44474
rect 21008 43722 21036 44746
rect 20996 43716 21048 43722
rect 20996 43658 21048 43664
rect 21008 42906 21036 43658
rect 20996 42900 21048 42906
rect 20996 42842 21048 42848
rect 21008 42634 21036 42842
rect 20996 42628 21048 42634
rect 20996 42570 21048 42576
rect 21100 41614 21128 51046
rect 21284 51046 21496 51074
rect 21284 44878 21312 51046
rect 21456 49088 21508 49094
rect 21456 49030 21508 49036
rect 21364 47456 21416 47462
rect 21364 47398 21416 47404
rect 21272 44872 21324 44878
rect 21270 44840 21272 44849
rect 21324 44840 21326 44849
rect 21270 44775 21326 44784
rect 21272 42764 21324 42770
rect 21272 42706 21324 42712
rect 21180 42560 21232 42566
rect 21180 42502 21232 42508
rect 21192 41682 21220 42502
rect 21284 42294 21312 42706
rect 21272 42288 21324 42294
rect 21272 42230 21324 42236
rect 21272 42152 21324 42158
rect 21272 42094 21324 42100
rect 21180 41676 21232 41682
rect 21180 41618 21232 41624
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 21088 41200 21140 41206
rect 21088 41142 21140 41148
rect 21100 40594 21128 41142
rect 21088 40588 21140 40594
rect 21088 40530 21140 40536
rect 21284 40458 21312 42094
rect 21376 40730 21404 47398
rect 21468 41274 21496 49030
rect 21560 44810 21588 53382
rect 21836 45558 21864 53926
rect 21928 53106 21956 56200
rect 22008 53440 22060 53446
rect 22008 53382 22060 53388
rect 21916 53100 21968 53106
rect 21916 53042 21968 53048
rect 22020 45966 22048 53382
rect 22296 53106 22324 56200
rect 22664 55214 22692 56200
rect 23032 56114 23060 56200
rect 23124 56114 23152 56222
rect 23032 56086 23152 56114
rect 22664 55186 22784 55214
rect 22756 54194 22784 55186
rect 22744 54188 22796 54194
rect 22744 54130 22796 54136
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53582 23336 56222
rect 24122 56200 24178 57000
rect 24490 56200 24546 57000
rect 24858 56200 24914 57000
rect 25226 56200 25282 57000
rect 25594 56200 25650 57000
rect 25962 56200 26018 57000
rect 24136 54262 24164 56200
rect 24124 54256 24176 54262
rect 24124 54198 24176 54204
rect 23756 54120 23808 54126
rect 23756 54062 23808 54068
rect 23388 53984 23440 53990
rect 23388 53926 23440 53932
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 23296 53440 23348 53446
rect 23296 53382 23348 53388
rect 22284 53100 22336 53106
rect 22284 53042 22336 53048
rect 22192 52896 22244 52902
rect 22192 52838 22244 52844
rect 22744 52896 22796 52902
rect 22744 52838 22796 52844
rect 22204 52601 22232 52838
rect 22190 52592 22246 52601
rect 22190 52527 22246 52536
rect 22468 46096 22520 46102
rect 22468 46038 22520 46044
rect 22100 46028 22152 46034
rect 22100 45970 22152 45976
rect 22008 45960 22060 45966
rect 22008 45902 22060 45908
rect 21824 45552 21876 45558
rect 21824 45494 21876 45500
rect 21916 44940 21968 44946
rect 21916 44882 21968 44888
rect 21548 44804 21600 44810
rect 21548 44746 21600 44752
rect 21560 44538 21588 44746
rect 21640 44736 21692 44742
rect 21640 44678 21692 44684
rect 21548 44532 21600 44538
rect 21548 44474 21600 44480
rect 21548 41472 21600 41478
rect 21548 41414 21600 41420
rect 21456 41268 21508 41274
rect 21456 41210 21508 41216
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21364 40724 21416 40730
rect 21364 40666 21416 40672
rect 21272 40452 21324 40458
rect 21272 40394 21324 40400
rect 21180 39976 21232 39982
rect 21180 39918 21232 39924
rect 21088 39500 21140 39506
rect 21088 39442 21140 39448
rect 21100 39030 21128 39442
rect 21088 39024 21140 39030
rect 21088 38966 21140 38972
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 21008 34678 21036 37606
rect 21100 37330 21128 38966
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 21192 37126 21220 39918
rect 21284 38418 21312 40394
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 21180 37120 21232 37126
rect 21180 37062 21232 37068
rect 21376 36768 21404 40666
rect 21468 40186 21496 40870
rect 21456 40180 21508 40186
rect 21456 40122 21508 40128
rect 21560 38350 21588 41414
rect 21652 39506 21680 44678
rect 21928 42158 21956 44882
rect 22008 44328 22060 44334
rect 22008 44270 22060 44276
rect 22020 43790 22048 44270
rect 22008 43784 22060 43790
rect 22008 43726 22060 43732
rect 22020 43246 22048 43726
rect 22008 43240 22060 43246
rect 22008 43182 22060 43188
rect 22020 42770 22048 43182
rect 22112 43110 22140 45970
rect 22376 45824 22428 45830
rect 22376 45766 22428 45772
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22296 43654 22324 44270
rect 22192 43648 22244 43654
rect 22192 43590 22244 43596
rect 22284 43648 22336 43654
rect 22284 43590 22336 43596
rect 22204 43450 22232 43590
rect 22192 43444 22244 43450
rect 22192 43386 22244 43392
rect 22100 43104 22152 43110
rect 22100 43046 22152 43052
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22008 42288 22060 42294
rect 22008 42230 22060 42236
rect 21916 42152 21968 42158
rect 21916 42094 21968 42100
rect 21916 42016 21968 42022
rect 21916 41958 21968 41964
rect 21732 41676 21784 41682
rect 21732 41618 21784 41624
rect 21640 39500 21692 39506
rect 21640 39442 21692 39448
rect 21548 38344 21600 38350
rect 21548 38286 21600 38292
rect 21456 38276 21508 38282
rect 21456 38218 21508 38224
rect 21192 36740 21404 36768
rect 21192 36106 21220 36740
rect 21364 36644 21416 36650
rect 21364 36586 21416 36592
rect 21272 36304 21324 36310
rect 21272 36246 21324 36252
rect 21180 36100 21232 36106
rect 21180 36042 21232 36048
rect 21088 35488 21140 35494
rect 21088 35430 21140 35436
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 21008 33114 21036 34138
rect 20996 33108 21048 33114
rect 20996 33050 21048 33056
rect 20996 32292 21048 32298
rect 20996 32234 21048 32240
rect 21008 31890 21036 32234
rect 21100 31890 21128 35430
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 21192 29714 21220 34682
rect 21284 32570 21312 36246
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21376 32502 21404 36586
rect 21468 36378 21496 38218
rect 21548 37664 21600 37670
rect 21548 37606 21600 37612
rect 21456 36372 21508 36378
rect 21456 36314 21508 36320
rect 21454 35728 21510 35737
rect 21454 35663 21510 35672
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21362 32056 21418 32065
rect 21362 31991 21364 32000
rect 21416 31991 21418 32000
rect 21364 31962 21416 31968
rect 21468 31872 21496 35663
rect 21560 35290 21588 37606
rect 21640 37324 21692 37330
rect 21640 37266 21692 37272
rect 21548 35284 21600 35290
rect 21548 35226 21600 35232
rect 21652 34474 21680 37266
rect 21744 36242 21772 41618
rect 21824 41608 21876 41614
rect 21822 41576 21824 41585
rect 21876 41576 21878 41585
rect 21822 41511 21878 41520
rect 21928 40050 21956 41958
rect 22020 41206 22048 42230
rect 22204 42158 22232 43386
rect 22192 42152 22244 42158
rect 22192 42094 22244 42100
rect 22008 41200 22060 41206
rect 22008 41142 22060 41148
rect 22100 41132 22152 41138
rect 22100 41074 22152 41080
rect 21916 40044 21968 40050
rect 21916 39986 21968 39992
rect 21824 39568 21876 39574
rect 21824 39510 21876 39516
rect 21836 39370 21864 39510
rect 21824 39364 21876 39370
rect 21824 39306 21876 39312
rect 21836 38214 21864 39306
rect 21916 39296 21968 39302
rect 21916 39238 21968 39244
rect 21824 38208 21876 38214
rect 21824 38150 21876 38156
rect 21836 37913 21864 38150
rect 21822 37904 21878 37913
rect 21822 37839 21878 37848
rect 21928 36378 21956 39238
rect 22008 38752 22060 38758
rect 22008 38694 22060 38700
rect 22020 36922 22048 38694
rect 22112 38486 22140 41074
rect 22204 39982 22232 42094
rect 22296 39982 22324 43590
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22284 39976 22336 39982
rect 22284 39918 22336 39924
rect 22192 39432 22244 39438
rect 22192 39374 22244 39380
rect 22100 38480 22152 38486
rect 22100 38422 22152 38428
rect 22204 37330 22232 39374
rect 22284 39296 22336 39302
rect 22284 39238 22336 39244
rect 22296 38554 22324 39238
rect 22388 39098 22416 45766
rect 22480 42362 22508 46038
rect 22652 43240 22704 43246
rect 22652 43182 22704 43188
rect 22560 42628 22612 42634
rect 22560 42570 22612 42576
rect 22468 42356 22520 42362
rect 22468 42298 22520 42304
rect 22572 41070 22600 42570
rect 22664 41426 22692 43182
rect 22756 41614 22784 52838
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23308 44946 23336 53382
rect 23296 44940 23348 44946
rect 23296 44882 23348 44888
rect 23400 44810 23428 53926
rect 23768 52698 23796 54062
rect 24872 53174 24900 56200
rect 25608 53650 25636 56200
rect 25596 53644 25648 53650
rect 25596 53586 25648 53592
rect 25872 53508 25924 53514
rect 25872 53450 25924 53456
rect 24860 53168 24912 53174
rect 24860 53110 24912 53116
rect 23756 52692 23808 52698
rect 23756 52634 23808 52640
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24124 51808 24176 51814
rect 24124 51750 24176 51756
rect 23480 44940 23532 44946
rect 23480 44882 23532 44888
rect 23388 44804 23440 44810
rect 23388 44746 23440 44752
rect 22836 44736 22888 44742
rect 22836 44678 22888 44684
rect 22744 41608 22796 41614
rect 22744 41550 22796 41556
rect 22664 41398 22784 41426
rect 22560 41064 22612 41070
rect 22560 41006 22612 41012
rect 22468 39364 22520 39370
rect 22468 39306 22520 39312
rect 22376 39092 22428 39098
rect 22376 39034 22428 39040
rect 22284 38548 22336 38554
rect 22284 38490 22336 38496
rect 22388 38010 22416 39034
rect 22480 38214 22508 39306
rect 22756 39030 22784 41398
rect 22848 41274 22876 44678
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 23204 41608 23256 41614
rect 23204 41550 23256 41556
rect 22836 41268 22888 41274
rect 22836 41210 22888 41216
rect 23216 41041 23244 41550
rect 23492 41206 23520 44882
rect 23848 44872 23900 44878
rect 23848 44814 23900 44820
rect 23860 44470 23888 44814
rect 23848 44464 23900 44470
rect 23848 44406 23900 44412
rect 23860 43722 23888 44406
rect 23848 43716 23900 43722
rect 23848 43658 23900 43664
rect 23860 43382 23888 43658
rect 23848 43376 23900 43382
rect 23848 43318 23900 43324
rect 23756 43240 23808 43246
rect 23756 43182 23808 43188
rect 23572 42560 23624 42566
rect 23572 42502 23624 42508
rect 23584 42294 23612 42502
rect 23572 42288 23624 42294
rect 23572 42230 23624 42236
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23202 41032 23258 41041
rect 23202 40967 23258 40976
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22836 40384 22888 40390
rect 22836 40326 22888 40332
rect 22848 39506 22876 40326
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22836 39500 22888 39506
rect 22836 39442 22888 39448
rect 22744 39024 22796 39030
rect 22744 38966 22796 38972
rect 22836 38956 22888 38962
rect 22836 38898 22888 38904
rect 22560 38548 22612 38554
rect 22560 38490 22612 38496
rect 22572 38418 22600 38490
rect 22560 38412 22612 38418
rect 22560 38354 22612 38360
rect 22468 38208 22520 38214
rect 22468 38150 22520 38156
rect 22572 38026 22600 38354
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22480 37998 22600 38026
rect 22744 38004 22796 38010
rect 22376 37460 22428 37466
rect 22376 37402 22428 37408
rect 22192 37324 22244 37330
rect 22192 37266 22244 37272
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 21732 36236 21784 36242
rect 21732 36178 21784 36184
rect 21640 34468 21692 34474
rect 21640 34410 21692 34416
rect 21744 33522 21772 36178
rect 22008 36100 22060 36106
rect 22008 36042 22060 36048
rect 22100 36100 22152 36106
rect 22100 36042 22152 36048
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21732 33516 21784 33522
rect 21732 33458 21784 33464
rect 21824 33108 21876 33114
rect 21824 33050 21876 33056
rect 21548 32768 21600 32774
rect 21548 32710 21600 32716
rect 21376 31844 21496 31872
rect 21376 30326 21404 31844
rect 21454 31784 21510 31793
rect 21454 31719 21456 31728
rect 21508 31719 21510 31728
rect 21456 31690 21508 31696
rect 21468 31210 21496 31690
rect 21456 31204 21508 31210
rect 21456 31146 21508 31152
rect 21364 30320 21416 30326
rect 21364 30262 21416 30268
rect 21272 29776 21324 29782
rect 21272 29718 21324 29724
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20904 25152 20956 25158
rect 20904 25094 20956 25100
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20548 21542 20668 21570
rect 20548 21078 20576 21542
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20640 20874 20760 20890
rect 20628 20868 20760 20874
rect 20680 20862 20760 20868
rect 20628 20810 20680 20816
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20456 16250 20484 18838
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20548 16046 20576 17478
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20088 15286 20208 15314
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19800 14000 19852 14006
rect 19800 13942 19852 13948
rect 19720 13824 19840 13852
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19352 12406 19472 12434
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19352 11830 19380 12242
rect 19444 12170 19472 12406
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19340 11824 19392 11830
rect 19392 11772 19472 11778
rect 19340 11766 19472 11772
rect 19352 11750 19472 11766
rect 19536 11762 19564 12650
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 19352 4622 19380 11562
rect 19444 11558 19472 11750
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 10674 19472 11494
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19628 5234 19656 12038
rect 19720 11218 19748 12582
rect 19812 11626 19840 13824
rect 20088 12374 20116 14214
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19996 11218 20024 11630
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19996 10810 20024 11154
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 5234 19748 6666
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 1170 18460 4014
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18340 1142 18460 1170
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 1142
rect 18524 898 18552 2314
rect 18432 870 18552 898
rect 18432 800 18460 870
rect 18800 800 18828 2790
rect 19168 800 19196 3402
rect 19444 3126 19472 5102
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19536 800 19564 5102
rect 19812 4486 19840 10610
rect 20088 6914 20116 12310
rect 20180 10062 20208 15286
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20272 13190 20300 13738
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20272 12918 20300 13126
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20364 11762 20392 15914
rect 20456 15570 20484 15914
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20640 14414 20668 20266
rect 20732 20262 20760 20862
rect 20824 20534 20852 25094
rect 20916 24274 20944 25094
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21008 21706 21036 29446
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 21100 26042 21128 29242
rect 21180 28620 21232 28626
rect 21284 28608 21312 29718
rect 21560 28778 21588 32710
rect 21732 31952 21784 31958
rect 21732 31894 21784 31900
rect 21744 30258 21772 31894
rect 21732 30252 21784 30258
rect 21732 30194 21784 30200
rect 21836 29730 21864 33050
rect 21928 32842 21956 33798
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 22020 32722 22048 36042
rect 22112 35154 22140 36042
rect 22100 35148 22152 35154
rect 22100 35090 22152 35096
rect 21928 32694 22048 32722
rect 21928 31822 21956 32694
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21744 29714 21864 29730
rect 21732 29708 21864 29714
rect 21784 29702 21864 29708
rect 21732 29650 21784 29656
rect 21560 28750 21772 28778
rect 21232 28580 21312 28608
rect 21180 28562 21232 28568
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 21100 24274 21128 25978
rect 21088 24268 21140 24274
rect 21192 24256 21220 28562
rect 21272 27056 21324 27062
rect 21272 26998 21324 27004
rect 21284 26246 21312 26998
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21284 25226 21312 26182
rect 21456 25764 21508 25770
rect 21456 25706 21508 25712
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21272 24268 21324 24274
rect 21192 24228 21272 24256
rect 21088 24210 21140 24216
rect 21272 24210 21324 24216
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20916 21678 21036 21706
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19990 20760 20198
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20916 18426 20944 21678
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20732 17270 20760 17546
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20732 14260 20760 17206
rect 20916 16522 20944 17274
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15434 20852 16050
rect 20916 16046 20944 16458
rect 21008 16182 21036 19450
rect 21100 19378 21128 23802
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20640 14232 20760 14260
rect 20640 13394 20668 14232
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20088 6886 20208 6914
rect 20180 5710 20208 6886
rect 20456 5846 20484 7686
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20548 4622 20576 13194
rect 20640 12918 20668 13330
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20640 12306 20668 12854
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20732 11218 20760 13670
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19904 800 19932 2858
rect 20272 800 20300 4014
rect 20364 2854 20392 4490
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20640 800 20668 5714
rect 20732 5710 20760 8842
rect 20824 7886 20852 14758
rect 20916 13326 20944 15982
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 21008 14074 21036 15574
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21100 13258 21128 15914
rect 21192 15026 21220 22918
rect 21284 22574 21312 24210
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21364 21548 21416 21554
rect 21364 21490 21416 21496
rect 21376 20874 21404 21490
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21376 17338 21404 18770
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21468 17218 21496 25706
rect 21652 25158 21680 26250
rect 21744 25838 21772 28750
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21732 25832 21784 25838
rect 21732 25774 21784 25780
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21560 21146 21588 21286
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21376 17190 21496 17218
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21284 13734 21312 14282
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21284 10674 21312 13466
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20824 6118 20852 7346
rect 20916 6458 20944 7346
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 21100 2922 21128 4490
rect 21284 3534 21312 7754
rect 21376 3602 21404 17190
rect 21652 16590 21680 20266
rect 21744 18766 21772 25638
rect 21928 23186 21956 27814
rect 22020 26042 22048 32166
rect 22112 28098 22140 35090
rect 22296 32570 22324 36722
rect 22388 36122 22416 37402
rect 22480 36582 22508 37998
rect 22744 37946 22796 37952
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 22664 37126 22692 37742
rect 22756 37466 22784 37946
rect 22744 37460 22796 37466
rect 22744 37402 22796 37408
rect 22848 37346 22876 38898
rect 23388 38888 23440 38894
rect 23388 38830 23440 38836
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 23296 38412 23348 38418
rect 23296 38354 23348 38360
rect 23308 37942 23336 38354
rect 23296 37936 23348 37942
rect 23296 37878 23348 37884
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22848 37318 22968 37346
rect 22940 37194 22968 37318
rect 22928 37188 22980 37194
rect 22928 37130 22980 37136
rect 22652 37120 22704 37126
rect 22652 37062 22704 37068
rect 23112 37120 23164 37126
rect 23112 37062 23164 37068
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22468 36576 22520 36582
rect 22468 36518 22520 36524
rect 22388 36094 22508 36122
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22190 32464 22246 32473
rect 22190 32399 22192 32408
rect 22244 32399 22246 32408
rect 22192 32370 22244 32376
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 22204 29646 22232 32166
rect 22388 32065 22416 35974
rect 22480 35154 22508 36094
rect 22572 35630 22600 36790
rect 22664 36718 22692 37062
rect 23124 36854 23152 37062
rect 23112 36848 23164 36854
rect 23112 36790 23164 36796
rect 22652 36712 22704 36718
rect 22652 36654 22704 36660
rect 22664 35630 22692 36654
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22848 36378 22876 36518
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22756 35698 22784 36314
rect 22836 36032 22888 36038
rect 22836 35974 22888 35980
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22652 35624 22704 35630
rect 22652 35566 22704 35572
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22468 34468 22520 34474
rect 22468 34410 22520 34416
rect 22480 33862 22508 34410
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22480 32978 22508 33798
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22572 32858 22600 34614
rect 22664 33454 22692 35566
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22652 33448 22704 33454
rect 22652 33390 22704 33396
rect 22480 32830 22600 32858
rect 22374 32056 22430 32065
rect 22374 31991 22430 32000
rect 22284 31952 22336 31958
rect 22480 31906 22508 32830
rect 22560 32768 22612 32774
rect 22560 32710 22612 32716
rect 22284 31894 22336 31900
rect 22296 30326 22324 31894
rect 22388 31878 22508 31906
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22388 29646 22416 31878
rect 22466 31784 22522 31793
rect 22466 31719 22522 31728
rect 22480 30666 22508 31719
rect 22468 30660 22520 30666
rect 22468 30602 22520 30608
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22376 29640 22428 29646
rect 22376 29582 22428 29588
rect 22192 28960 22244 28966
rect 22192 28902 22244 28908
rect 22204 28558 22232 28902
rect 22192 28552 22244 28558
rect 22192 28494 22244 28500
rect 22112 28070 22324 28098
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 22112 26194 22140 27882
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22204 27130 22232 27406
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 22204 26926 22232 27066
rect 22192 26920 22244 26926
rect 22192 26862 22244 26868
rect 22204 26450 22232 26862
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22112 26166 22232 26194
rect 22098 26072 22154 26081
rect 22008 26036 22060 26042
rect 22098 26007 22154 26016
rect 22008 25978 22060 25984
rect 22112 25702 22140 26007
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 22112 23118 22140 24550
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 13870 21496 15846
rect 21836 15570 21864 19722
rect 21928 16522 21956 19994
rect 22112 19378 22140 22918
rect 22204 22642 22232 26166
rect 22296 26042 22324 28070
rect 22480 27554 22508 29786
rect 22572 28218 22600 32710
rect 22664 30802 22692 33390
rect 22756 31906 22784 35430
rect 22848 32230 22876 35974
rect 23308 35494 23336 37878
rect 23400 37806 23428 38830
rect 23492 38554 23520 41142
rect 23584 40594 23612 42230
rect 23664 40928 23716 40934
rect 23664 40870 23716 40876
rect 23572 40588 23624 40594
rect 23572 40530 23624 40536
rect 23676 40526 23704 40870
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23572 40384 23624 40390
rect 23572 40326 23624 40332
rect 23664 40384 23716 40390
rect 23664 40326 23716 40332
rect 23480 38548 23532 38554
rect 23480 38490 23532 38496
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23308 35154 23336 35430
rect 23204 35148 23256 35154
rect 23204 35090 23256 35096
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 23216 35034 23244 35090
rect 23216 35006 23336 35034
rect 23204 34944 23256 34950
rect 23204 34886 23256 34892
rect 23216 34610 23244 34886
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23308 34218 23336 35006
rect 23400 34746 23428 37062
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 36242 23520 36518
rect 23480 36236 23532 36242
rect 23480 36178 23532 36184
rect 23492 35766 23520 36178
rect 23480 35760 23532 35766
rect 23480 35702 23532 35708
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23308 34190 23428 34218
rect 23296 34128 23348 34134
rect 23296 34070 23348 34076
rect 23308 33590 23336 34070
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23020 33108 23072 33114
rect 23020 33050 23072 33056
rect 23032 32842 23060 33050
rect 23112 32972 23164 32978
rect 23112 32914 23164 32920
rect 23124 32858 23152 32914
rect 23308 32910 23336 33526
rect 23400 33114 23428 34190
rect 23584 34066 23612 40326
rect 23676 39642 23704 40326
rect 23664 39636 23716 39642
rect 23664 39578 23716 39584
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23676 36242 23704 38150
rect 23768 38010 23796 43182
rect 23860 42906 23888 43318
rect 23848 42900 23900 42906
rect 23848 42842 23900 42848
rect 23860 42634 23888 42842
rect 23848 42628 23900 42634
rect 23848 42570 23900 42576
rect 23940 41608 23992 41614
rect 23940 41550 23992 41556
rect 23848 40180 23900 40186
rect 23848 40122 23900 40128
rect 23756 38004 23808 38010
rect 23756 37946 23808 37952
rect 23754 37632 23810 37641
rect 23754 37567 23810 37576
rect 23768 37262 23796 37567
rect 23756 37256 23808 37262
rect 23756 37198 23808 37204
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 23664 36236 23716 36242
rect 23664 36178 23716 36184
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35290 23704 35974
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23388 32972 23440 32978
rect 23388 32914 23440 32920
rect 23296 32904 23348 32910
rect 23020 32836 23072 32842
rect 23124 32830 23244 32858
rect 23296 32846 23348 32852
rect 23020 32778 23072 32784
rect 23216 32366 23244 32830
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23204 32360 23256 32366
rect 23204 32302 23256 32308
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31958 23336 32370
rect 23296 31952 23348 31958
rect 22926 31920 22982 31929
rect 22756 31878 22876 31906
rect 22848 31346 22876 31878
rect 23296 31894 23348 31900
rect 22926 31855 22982 31864
rect 23020 31884 23072 31890
rect 22940 31686 22968 31855
rect 23020 31826 23072 31832
rect 23032 31793 23060 31826
rect 23018 31784 23074 31793
rect 23018 31719 23074 31728
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22940 31226 22968 31622
rect 22848 31198 22968 31226
rect 22652 30796 22704 30802
rect 22652 30738 22704 30744
rect 22664 30258 22692 30738
rect 22652 30252 22704 30258
rect 22652 30194 22704 30200
rect 22652 30116 22704 30122
rect 22652 30058 22704 30064
rect 22664 28626 22692 30058
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22560 28212 22612 28218
rect 22560 28154 22612 28160
rect 22480 27526 22600 27554
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22480 27130 22508 27338
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22468 26920 22520 26926
rect 22468 26862 22520 26868
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22296 25401 22324 25842
rect 22282 25392 22338 25401
rect 22282 25327 22338 25336
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22204 20942 22232 21422
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22204 19281 22232 19382
rect 22190 19272 22246 19281
rect 22190 19207 22246 19216
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 18222 22048 18702
rect 22112 18290 22140 19110
rect 22192 18896 22244 18902
rect 22192 18838 22244 18844
rect 22204 18290 22232 18838
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 22020 17202 22048 18158
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 22112 15570 22140 16934
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22204 15026 22232 18022
rect 22296 17678 22324 25162
rect 22388 24750 22416 26522
rect 22480 24954 22508 26862
rect 22572 25242 22600 27526
rect 22664 25362 22692 28358
rect 22848 28082 22876 31198
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23308 28762 23336 29446
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22848 26568 22876 28018
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23308 27674 23336 27814
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23400 27554 23428 32914
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23492 31890 23520 32166
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 23492 29714 23520 29990
rect 23480 29708 23532 29714
rect 23480 29650 23532 29656
rect 23584 29578 23612 32710
rect 23572 29572 23624 29578
rect 23572 29514 23624 29520
rect 23676 28150 23704 33798
rect 23768 33590 23796 36314
rect 23860 33998 23888 40122
rect 23952 35737 23980 41550
rect 24030 40352 24086 40361
rect 24030 40287 24086 40296
rect 24044 39438 24072 40287
rect 24032 39432 24084 39438
rect 24032 39374 24084 39380
rect 24136 36106 24164 51750
rect 24504 44878 24532 52430
rect 25136 52012 25188 52018
rect 25136 51954 25188 51960
rect 25148 51921 25176 51954
rect 25134 51912 25190 51921
rect 25134 51847 25190 51856
rect 25044 51400 25096 51406
rect 25044 51342 25096 51348
rect 25056 51241 25084 51342
rect 25596 51264 25648 51270
rect 25042 51232 25098 51241
rect 25596 51206 25648 51212
rect 25042 51167 25098 51176
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25044 50312 25096 50318
rect 25044 50254 25096 50260
rect 25056 49881 25084 50254
rect 25042 49872 25098 49881
rect 25042 49807 25098 49816
rect 25044 49224 25096 49230
rect 25042 49192 25044 49201
rect 25096 49192 25098 49201
rect 25042 49127 25098 49136
rect 25044 48748 25096 48754
rect 25044 48690 25096 48696
rect 25056 48521 25084 48690
rect 25136 48544 25188 48550
rect 25042 48512 25098 48521
rect 25136 48486 25188 48492
rect 25042 48447 25098 48456
rect 25044 48136 25096 48142
rect 25044 48078 25096 48084
rect 25056 47841 25084 48078
rect 25042 47832 25098 47841
rect 25042 47767 25098 47776
rect 25044 47660 25096 47666
rect 25044 47602 25096 47608
rect 25056 47161 25084 47602
rect 25042 47152 25098 47161
rect 25042 47087 25098 47096
rect 24676 45960 24728 45966
rect 24676 45902 24728 45908
rect 24584 45484 24636 45490
rect 24584 45426 24636 45432
rect 24596 45082 24624 45426
rect 24688 45121 24716 45902
rect 24766 45792 24822 45801
rect 24766 45727 24822 45736
rect 24780 45422 24808 45727
rect 24768 45416 24820 45422
rect 24768 45358 24820 45364
rect 24674 45112 24730 45121
rect 24584 45076 24636 45082
rect 24674 45047 24730 45056
rect 24584 45018 24636 45024
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 24858 44432 24914 44441
rect 24858 44367 24860 44376
rect 24912 44367 24914 44376
rect 24860 44338 24912 44344
rect 24952 44192 25004 44198
rect 24952 44134 25004 44140
rect 24768 43784 24820 43790
rect 24768 43726 24820 43732
rect 24584 42628 24636 42634
rect 24584 42570 24636 42576
rect 24596 42294 24624 42570
rect 24780 42401 24808 43726
rect 24860 43308 24912 43314
rect 24860 43250 24912 43256
rect 24872 43081 24900 43250
rect 24858 43072 24914 43081
rect 24858 43007 24914 43016
rect 24766 42392 24822 42401
rect 24766 42327 24822 42336
rect 24584 42288 24636 42294
rect 24584 42230 24636 42236
rect 24596 41562 24624 42230
rect 24964 41750 24992 44134
rect 25148 43858 25176 48486
rect 25412 48000 25464 48006
rect 25412 47942 25464 47948
rect 25320 44396 25372 44402
rect 25320 44338 25372 44344
rect 25136 43852 25188 43858
rect 25136 43794 25188 43800
rect 25332 43761 25360 44338
rect 25318 43752 25374 43761
rect 25318 43687 25374 43696
rect 25320 42696 25372 42702
rect 25320 42638 25372 42644
rect 25228 42560 25280 42566
rect 25228 42502 25280 42508
rect 24952 41744 25004 41750
rect 24952 41686 25004 41692
rect 24504 41534 24624 41562
rect 24504 41206 24532 41534
rect 24492 41200 24544 41206
rect 24412 41160 24492 41188
rect 24412 40458 24440 41160
rect 24492 41142 24544 41148
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 24952 40520 25004 40526
rect 24952 40462 25004 40468
rect 24400 40452 24452 40458
rect 24400 40394 24452 40400
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24216 38888 24268 38894
rect 24216 38830 24268 38836
rect 24228 38010 24256 38830
rect 24216 38004 24268 38010
rect 24216 37946 24268 37952
rect 24228 36242 24256 37946
rect 24216 36236 24268 36242
rect 24216 36178 24268 36184
rect 24124 36100 24176 36106
rect 24124 36042 24176 36048
rect 23938 35728 23994 35737
rect 23938 35663 23994 35672
rect 24320 34678 24348 39238
rect 24412 39030 24440 40394
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 24872 39681 24900 39986
rect 24858 39672 24914 39681
rect 24858 39607 24914 39616
rect 24964 39438 24992 40462
rect 25056 39506 25084 40870
rect 25136 39908 25188 39914
rect 25136 39850 25188 39856
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 24952 39432 25004 39438
rect 24952 39374 25004 39380
rect 25044 39296 25096 39302
rect 25044 39238 25096 39244
rect 24400 39024 24452 39030
rect 24452 38972 24532 38978
rect 24400 38966 24532 38972
rect 24412 38950 24532 38966
rect 24504 37942 24532 38950
rect 24492 37936 24544 37942
rect 24492 37878 24544 37884
rect 24504 37194 24532 37878
rect 24860 37256 24912 37262
rect 24860 37198 24912 37204
rect 24492 37188 24544 37194
rect 24492 37130 24544 37136
rect 24504 36854 24532 37130
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 24596 36922 24624 37062
rect 24872 36961 24900 37198
rect 24858 36952 24914 36961
rect 24584 36916 24636 36922
rect 24858 36887 24914 36896
rect 24584 36858 24636 36864
rect 24492 36848 24544 36854
rect 24492 36790 24544 36796
rect 24504 35766 24532 36790
rect 24860 36576 24912 36582
rect 24860 36518 24912 36524
rect 24492 35760 24544 35766
rect 24492 35702 24544 35708
rect 24308 34672 24360 34678
rect 24308 34614 24360 34620
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 24504 33930 24532 35702
rect 24872 34134 24900 36518
rect 25056 36174 25084 39238
rect 25148 39001 25176 39850
rect 25134 38992 25190 39001
rect 25134 38927 25190 38936
rect 25136 38208 25188 38214
rect 25136 38150 25188 38156
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 25148 35086 25176 38150
rect 25240 37670 25268 42502
rect 25332 41721 25360 42638
rect 25318 41712 25374 41721
rect 25318 41647 25374 41656
rect 25320 41608 25372 41614
rect 25320 41550 25372 41556
rect 25332 38321 25360 41550
rect 25424 39370 25452 47942
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25412 39364 25464 39370
rect 25412 39306 25464 39312
rect 25412 38344 25464 38350
rect 25318 38312 25374 38321
rect 25412 38286 25464 38292
rect 25318 38247 25374 38256
rect 25228 37664 25280 37670
rect 25228 37606 25280 37612
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25332 35601 25360 36722
rect 25424 36281 25452 38286
rect 25516 36718 25544 43590
rect 25504 36712 25556 36718
rect 25504 36654 25556 36660
rect 25410 36272 25466 36281
rect 25410 36207 25466 36216
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25318 35592 25374 35601
rect 25318 35527 25374 35536
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 24860 34128 24912 34134
rect 24860 34070 24912 34076
rect 24492 33924 24544 33930
rect 24492 33866 24544 33872
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 23756 33584 23808 33590
rect 23756 33526 23808 33532
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23768 30054 23796 33390
rect 23860 31226 23888 33594
rect 24504 33590 24532 33866
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24308 32224 24360 32230
rect 24308 32166 24360 32172
rect 24032 31816 24084 31822
rect 24032 31758 24084 31764
rect 24044 31521 24072 31758
rect 24030 31512 24086 31521
rect 24030 31447 24086 31456
rect 23860 31198 23980 31226
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 29714 23796 29990
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23308 27538 23428 27554
rect 23296 27532 23428 27538
rect 23348 27526 23428 27532
rect 23296 27474 23348 27480
rect 23308 26874 23336 27474
rect 23216 26846 23336 26874
rect 23216 26790 23244 26846
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23308 26586 23336 26846
rect 23492 26761 23520 28018
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23768 27606 23796 27950
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 23572 26784 23624 26790
rect 23478 26752 23534 26761
rect 23572 26726 23624 26732
rect 23478 26687 23534 26696
rect 23296 26580 23348 26586
rect 22848 26540 22968 26568
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22756 26330 22784 26386
rect 22756 26302 22876 26330
rect 22744 25696 22796 25702
rect 22744 25638 22796 25644
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22572 25214 22692 25242
rect 22664 25158 22692 25214
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22376 24744 22428 24750
rect 22376 24686 22428 24692
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 23186 22416 24550
rect 22480 24410 22508 24754
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22388 21146 22416 22714
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22388 19174 22416 20878
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22480 18358 22508 22374
rect 22572 20534 22600 25094
rect 22756 23338 22784 25638
rect 22848 24750 22876 26302
rect 22940 26081 22968 26540
rect 23296 26522 23348 26528
rect 22926 26072 22982 26081
rect 22926 26007 22982 26016
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22664 23310 22784 23338
rect 22664 22982 22692 23310
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22664 22166 22692 22510
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22664 21554 22692 22102
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22664 20466 22692 21490
rect 22756 20942 22784 23190
rect 22848 22574 22876 24686
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22664 19990 22692 20402
rect 22848 20262 22876 21558
rect 22940 21486 22968 22170
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22940 20602 22968 20742
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22296 13938 22324 15642
rect 22388 14414 22416 18226
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22480 14958 22508 18090
rect 22572 16182 22600 18770
rect 23308 18630 23336 25774
rect 23480 25764 23532 25770
rect 23480 25706 23532 25712
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 23400 23746 23428 25298
rect 23492 23866 23520 25706
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23400 23718 23520 23746
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 23400 23361 23428 23598
rect 23386 23352 23442 23361
rect 23386 23287 23442 23296
rect 23492 22778 23520 23718
rect 23584 23118 23612 26726
rect 23768 24834 23796 27542
rect 23860 27470 23888 31078
rect 23952 28762 23980 31198
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 24044 30190 24072 30534
rect 24228 30326 24256 30738
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24032 30184 24084 30190
rect 24032 30126 24084 30132
rect 24032 29776 24084 29782
rect 24032 29718 24084 29724
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 24044 28082 24072 29718
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24136 28801 24164 29106
rect 24122 28792 24178 28801
rect 24122 28727 24178 28736
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 24228 27962 24256 30262
rect 24136 27934 24256 27962
rect 23940 27872 23992 27878
rect 23940 27814 23992 27820
rect 23848 27464 23900 27470
rect 23848 27406 23900 27412
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23860 26586 23888 27270
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23952 25294 23980 27814
rect 24136 27402 24164 27934
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 24136 27062 24164 27338
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 24136 26314 24164 26998
rect 24124 26308 24176 26314
rect 24044 26268 24124 26296
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 24044 24886 24072 26268
rect 24124 26250 24176 26256
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 23676 24806 23796 24834
rect 24032 24880 24084 24886
rect 24032 24822 24084 24828
rect 23676 24750 23704 24806
rect 23664 24744 23716 24750
rect 23664 24686 23716 24692
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23492 21010 23520 22714
rect 24044 22710 24072 24822
rect 24136 23730 24164 25094
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 24044 22094 24072 22646
rect 23768 22066 24072 22094
rect 23768 21690 23796 22066
rect 24228 22030 24256 27814
rect 24320 26314 24348 32166
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24412 30569 24440 31282
rect 24504 30802 24532 33526
rect 24492 30796 24544 30802
rect 24492 30738 24544 30744
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 24398 30560 24454 30569
rect 24398 30495 24454 30504
rect 24504 30433 24532 30602
rect 24490 30424 24546 30433
rect 24490 30359 24546 30368
rect 24596 29238 24624 33798
rect 24860 32904 24912 32910
rect 24858 32872 24860 32881
rect 24912 32872 24914 32881
rect 24858 32807 24914 32816
rect 24676 31952 24728 31958
rect 24676 31894 24728 31900
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24308 26308 24360 26314
rect 24308 26250 24360 26256
rect 24412 24206 24440 28970
rect 24688 27062 24716 31894
rect 25056 30394 25084 34682
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 33561 25360 34546
rect 25424 34241 25452 35022
rect 25516 34921 25544 36110
rect 25502 34912 25558 34921
rect 25502 34847 25558 34856
rect 25410 34232 25466 34241
rect 25410 34167 25466 34176
rect 25318 33552 25374 33561
rect 25318 33487 25374 33496
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25136 32768 25188 32774
rect 25134 32736 25136 32745
rect 25188 32736 25190 32745
rect 25134 32671 25190 32680
rect 25136 32564 25188 32570
rect 25136 32506 25188 32512
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25148 29850 25176 32506
rect 25332 32201 25360 32846
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25318 32192 25374 32201
rect 25318 32127 25374 32136
rect 25228 31204 25280 31210
rect 25228 31146 25280 31152
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 24860 28552 24912 28558
rect 24860 28494 24912 28500
rect 24872 28121 24900 28494
rect 24858 28112 24914 28121
rect 24858 28047 24914 28056
rect 24950 27432 25006 27441
rect 24860 27396 24912 27402
rect 24950 27367 25006 27376
rect 24860 27338 24912 27344
rect 24676 27056 24728 27062
rect 24676 26998 24728 27004
rect 24766 26072 24822 26081
rect 24766 26007 24822 26016
rect 24780 24206 24808 26007
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24872 23798 24900 27338
rect 24964 26382 24992 27367
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24964 24041 24992 24074
rect 24950 24032 25006 24041
rect 24950 23967 25006 23976
rect 24860 23792 24912 23798
rect 24860 23734 24912 23740
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24950 21992 25006 22001
rect 24950 21927 24952 21936
rect 25004 21927 25006 21936
rect 24952 21898 25004 21904
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23492 20602 23520 20946
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23768 20534 23796 21626
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24674 21312 24730 21321
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 22664 18154 22692 18566
rect 23308 18426 23336 18566
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22652 18148 22704 18154
rect 22652 18090 22704 18096
rect 22756 16998 22784 18294
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17921 23428 18022
rect 23386 17912 23442 17921
rect 23386 17847 23442 17856
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22848 16810 22876 17070
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22756 16782 22876 16810
rect 22756 16182 22784 16782
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21008 800 21036 2790
rect 21468 2446 21496 13670
rect 21560 4214 21588 13874
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21652 13258 21680 13330
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22112 12442 22140 12786
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22388 11898 22416 12174
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22572 11354 22600 11698
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22204 9586 22232 11222
rect 22664 11218 22692 13670
rect 22848 12850 22876 16594
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 13530 23336 13942
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22756 9042 22784 10950
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22848 8922 22876 11562
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22756 8894 22876 8922
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21548 4208 21600 4214
rect 21548 4150 21600 4156
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21560 2122 21588 3946
rect 21376 2094 21588 2122
rect 21376 800 21404 2094
rect 21744 800 21772 5578
rect 22020 3398 22048 6666
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22112 5914 22140 6258
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22204 3210 22232 6190
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22112 3182 22232 3210
rect 22112 800 22140 3182
rect 22296 2854 22324 5102
rect 22388 4321 22416 6326
rect 22374 4312 22430 4321
rect 22374 4247 22430 4256
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22480 800 22508 7278
rect 22756 5574 22784 8894
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 6798 22876 8774
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23308 7886 23336 11290
rect 23400 11082 23428 14214
rect 23492 13938 23520 19178
rect 23768 18698 23796 20470
rect 24596 18766 24624 21286
rect 24674 21247 24730 21256
rect 24688 19310 24716 21247
rect 24950 20632 25006 20641
rect 24950 20567 25006 20576
rect 24858 19952 24914 19961
rect 24964 19922 24992 20567
rect 24858 19887 24914 19896
rect 24952 19916 25004 19922
rect 24872 19446 24900 19887
rect 24952 19858 25004 19864
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 25056 19378 25084 26250
rect 25240 25974 25268 31146
rect 25424 30841 25452 32370
rect 25608 31754 25636 51206
rect 25688 50720 25740 50726
rect 25688 50662 25740 50668
rect 25700 38486 25728 50662
rect 25780 50176 25832 50182
rect 25780 50118 25832 50124
rect 25792 39574 25820 50118
rect 25780 39568 25832 39574
rect 25780 39510 25832 39516
rect 25688 38480 25740 38486
rect 25688 38422 25740 38428
rect 25596 31748 25648 31754
rect 25596 31690 25648 31696
rect 25884 31414 25912 53450
rect 25964 53100 26016 53106
rect 25964 53042 26016 53048
rect 25872 31408 25924 31414
rect 25872 31350 25924 31356
rect 25976 30870 26004 53042
rect 25964 30864 26016 30870
rect 25410 30832 25466 30841
rect 25964 30806 26016 30812
rect 25410 30767 25466 30776
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25318 29472 25374 29481
rect 25318 29407 25374 29416
rect 25332 28558 25360 29407
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25228 25968 25280 25974
rect 25228 25910 25280 25916
rect 25228 25764 25280 25770
rect 25228 25706 25280 25712
rect 25134 24712 25190 24721
rect 25134 24647 25190 24656
rect 25148 23798 25176 24647
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25240 19854 25268 25706
rect 26056 23044 26108 23050
rect 26056 22986 26108 22992
rect 26068 22681 26096 22986
rect 26054 22672 26110 22681
rect 26054 22607 26110 22616
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 23756 18692 23808 18698
rect 23756 18634 23808 18640
rect 23768 18358 23796 18634
rect 24216 18624 24268 18630
rect 23846 18592 23902 18601
rect 24216 18566 24268 18572
rect 23846 18527 23902 18536
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23768 17270 23796 18294
rect 23860 17746 23888 18527
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23756 17264 23808 17270
rect 23756 17206 23808 17212
rect 23846 17232 23902 17241
rect 23846 17167 23902 17176
rect 23860 16590 23888 17167
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23768 10130 23796 13126
rect 23860 11762 23888 16186
rect 23940 15632 23992 15638
rect 23940 15574 23992 15580
rect 23952 13326 23980 15574
rect 24228 15026 24256 18566
rect 24766 16552 24822 16561
rect 24766 16487 24822 16496
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15434 24440 15846
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24780 14958 24808 16487
rect 24858 15872 24914 15881
rect 24858 15807 24914 15816
rect 24872 15570 24900 15807
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 25134 15192 25190 15201
rect 25134 15127 25190 15136
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24872 14521 24900 15030
rect 24858 14512 24914 14521
rect 24858 14447 24914 14456
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24596 12238 24624 14010
rect 25148 14006 25176 15127
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24674 13152 24730 13161
rect 24674 13087 24730 13096
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23492 3602 23520 6666
rect 23584 5030 23612 9522
rect 23860 8498 23888 10950
rect 23952 10674 23980 11494
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24596 10062 24624 12038
rect 24688 11694 24716 13087
rect 24780 12782 24808 13767
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24872 12481 24900 12854
rect 24858 12472 24914 12481
rect 24858 12407 24914 12416
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 25332 11801 25360 12106
rect 25318 11792 25374 11801
rect 25318 11727 25374 11736
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24766 11112 24822 11121
rect 24766 11047 24822 11056
rect 24780 10606 24808 11047
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24766 10432 24822 10441
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 24044 8974 24072 9318
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 24136 6322 24164 8774
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24504 6914 24532 8366
rect 24596 7410 24624 9862
rect 24688 7886 24716 10406
rect 24766 10367 24822 10376
rect 24780 9518 24808 10367
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 24964 9761 24992 9930
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 25134 9072 25190 9081
rect 25134 9007 25190 9016
rect 25148 8566 25176 9007
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24766 8392 24822 8401
rect 24766 8327 24822 8336
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24504 6886 24624 6914
rect 24490 6760 24546 6769
rect 24490 6695 24492 6704
rect 24544 6695 24546 6704
rect 24492 6666 24544 6672
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24490 5672 24546 5681
rect 24490 5607 24492 5616
rect 24544 5607 24546 5616
rect 24492 5578 24544 5584
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 800 22876 3334
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2530 23336 3538
rect 23768 3194 23796 4558
rect 23860 4146 23888 5510
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23216 2502 23336 2530
rect 23216 800 23244 2502
rect 23584 800 23612 2994
rect 23952 800 23980 3062
rect 24320 800 24348 3402
rect 24504 2990 24532 5578
rect 24596 3482 24624 6886
rect 24688 5234 24716 7686
rect 24780 7342 24808 8327
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24766 7032 24822 7041
rect 24766 6967 24822 6976
rect 24780 6254 24808 6967
rect 24872 6866 24900 8502
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7721 24992 7754
rect 24950 7712 25006 7721
rect 24950 7647 25006 7656
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6361 24992 6734
rect 24950 6352 25006 6361
rect 24950 6287 25006 6296
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 5914 24808 6054
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 24766 5672 24822 5681
rect 24766 5607 24822 5616
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24780 5166 24808 5607
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 25318 4992 25374 5001
rect 25318 4927 25374 4936
rect 25332 4826 25360 4927
rect 25320 4820 25372 4826
rect 25320 4762 25372 4768
rect 24596 3454 24716 3482
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24688 800 24716 3454
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 25056 800 25084 2858
rect 25424 800 25452 7414
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
<< via2 >>
rect 938 50360 994 50416
rect 1306 52672 1362 52728
rect 2778 54984 2834 55040
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 938 48068 994 48104
rect 938 48048 940 48068
rect 940 48048 992 48068
rect 992 48048 994 48068
rect 938 45736 994 45792
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 1674 41112 1730 41168
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 938 38800 994 38856
rect 938 36488 994 36544
rect 1766 34176 1822 34232
rect 938 31864 994 31920
rect 1306 29552 1362 29608
rect 1306 27240 1362 27296
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 1306 24928 1362 24984
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 1306 22616 1362 22672
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 1306 20340 1308 20360
rect 1308 20340 1360 20360
rect 1360 20340 1362 20360
rect 1306 20304 1362 20340
rect 1306 17992 1362 18048
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 1306 15680 1362 15736
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2778 13368 2834 13424
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2778 11056 2834 11112
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3054 8744 3110 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3146 6432 3202 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3238 4120 3294 4176
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2778 1808 2834 1864
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7194 44240 7250 44296
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 5078 2896 5134 2952
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 10230 42880 10286 42936
rect 9034 36080 9090 36136
rect 9034 31864 9090 31920
rect 10322 41384 10378 41440
rect 9402 31864 9458 31920
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7838 5616 7894 5672
rect 7654 4120 7710 4176
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 8390 3732 8446 3768
rect 8390 3712 8392 3732
rect 8392 3712 8444 3732
rect 8444 3712 8446 3732
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 10046 27240 10102 27296
rect 10874 34584 10930 34640
rect 10414 21428 10416 21448
rect 10416 21428 10468 21448
rect 10468 21428 10470 21448
rect 10414 21392 10470 21428
rect 11794 44240 11850 44296
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 14830 53932 14832 53952
rect 14832 53932 14884 53952
rect 14884 53932 14886 53952
rect 14830 53896 14886 53932
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 11886 35944 11942 36000
rect 11886 33768 11942 33824
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12070 27920 12126 27976
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12714 31628 12716 31648
rect 12716 31628 12768 31648
rect 12768 31628 12770 31648
rect 12714 31592 12770 31628
rect 12254 27376 12310 27432
rect 12070 24948 12126 24984
rect 12070 24928 12072 24948
rect 12072 24928 12124 24948
rect 12124 24928 12126 24948
rect 12438 25200 12494 25256
rect 12070 21936 12126 21992
rect 12346 21836 12348 21856
rect 12348 21836 12400 21856
rect 12400 21836 12402 21856
rect 12346 21800 12402 21836
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 13634 35148 13690 35184
rect 13634 35128 13636 35148
rect 13636 35128 13688 35148
rect 13688 35128 13690 35148
rect 13358 30540 13360 30560
rect 13360 30540 13412 30560
rect 13412 30540 13414 30560
rect 13358 30504 13414 30540
rect 12990 30096 13046 30152
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 13174 27276 13176 27296
rect 13176 27276 13228 27296
rect 13228 27276 13230 27296
rect 13174 27240 13230 27276
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12806 25200 12862 25256
rect 12898 25064 12954 25120
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12898 22480 12954 22536
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12346 18400 12402 18456
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 13450 21428 13452 21448
rect 13452 21428 13504 21448
rect 13504 21428 13506 21448
rect 13450 21392 13506 21428
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 14554 52536 14610 52592
rect 15566 46008 15622 46064
rect 14278 32000 14334 32056
rect 13910 21564 13912 21584
rect 13912 21564 13964 21584
rect 13964 21564 13966 21584
rect 13910 21528 13966 21564
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 14002 16224 14058 16280
rect 15290 37712 15346 37768
rect 15290 36216 15346 36272
rect 15290 30132 15292 30152
rect 15292 30132 15344 30152
rect 15344 30132 15346 30152
rect 15290 30096 15346 30132
rect 15106 26868 15108 26888
rect 15108 26868 15160 26888
rect 15160 26868 15162 26888
rect 15106 26832 15162 26868
rect 14554 21392 14610 21448
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 16210 38156 16212 38176
rect 16212 38156 16264 38176
rect 16264 38156 16266 38176
rect 16210 38120 16266 38156
rect 16210 36660 16212 36680
rect 16212 36660 16264 36680
rect 16264 36660 16266 36680
rect 16210 36624 16266 36660
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 18418 46416 18474 46472
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 16946 37712 17002 37768
rect 16762 32444 16764 32464
rect 16764 32444 16816 32464
rect 16816 32444 16818 32464
rect 16762 32408 16818 32444
rect 16486 29008 16542 29064
rect 16026 27276 16028 27296
rect 16028 27276 16080 27296
rect 16080 27276 16082 27296
rect 16026 27240 16082 27276
rect 15566 21800 15622 21856
rect 15382 16496 15438 16552
rect 15198 16224 15254 16280
rect 16118 21664 16174 21720
rect 17038 32136 17094 32192
rect 17314 32564 17370 32600
rect 17314 32544 17316 32564
rect 17316 32544 17368 32564
rect 17368 32544 17370 32564
rect 17590 37068 17592 37088
rect 17592 37068 17644 37088
rect 17644 37068 17646 37088
rect 17590 37032 17646 37068
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17590 36488 17646 36544
rect 17682 36352 17738 36408
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17866 37748 17868 37768
rect 17868 37748 17920 37768
rect 17920 37748 17922 37768
rect 17866 37712 17922 37748
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 18326 36624 18382 36680
rect 18510 36660 18512 36680
rect 18512 36660 18564 36680
rect 18564 36660 18566 36680
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 18510 36624 18566 36660
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17682 32136 17738 32192
rect 17590 29452 17592 29472
rect 17592 29452 17644 29472
rect 17644 29452 17646 29472
rect 17590 29416 17646 29452
rect 16670 24792 16726 24848
rect 16946 22208 17002 22264
rect 17130 22208 17186 22264
rect 17038 19388 17040 19408
rect 17040 19388 17092 19408
rect 17092 19388 17094 19408
rect 17038 19352 17094 19388
rect 17314 20576 17370 20632
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17958 27512 18014 27568
rect 17866 27376 17922 27432
rect 19798 45772 19800 45792
rect 19800 45772 19852 45792
rect 19852 45772 19854 45792
rect 18878 36624 18934 36680
rect 18602 35672 18658 35728
rect 19154 40024 19210 40080
rect 18418 27956 18420 27976
rect 18420 27956 18472 27976
rect 18472 27956 18474 27976
rect 18418 27920 18474 27956
rect 18418 27532 18474 27568
rect 18418 27512 18420 27532
rect 18420 27512 18472 27532
rect 18472 27512 18474 27532
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17590 23432 17646 23488
rect 17498 22072 17554 22128
rect 17222 20440 17278 20496
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17866 21936 17922 21992
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 19798 45736 19854 45772
rect 20626 45600 20682 45656
rect 18970 29280 19026 29336
rect 19154 30252 19210 30288
rect 19154 30232 19156 30252
rect 19156 30232 19208 30252
rect 19208 30232 19210 30252
rect 18878 27920 18934 27976
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18786 19352 18842 19408
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 19522 34584 19578 34640
rect 19522 29300 19578 29336
rect 19522 29280 19524 29300
rect 19524 29280 19576 29300
rect 19576 29280 19578 29300
rect 20442 36216 20498 36272
rect 20350 36100 20406 36136
rect 20350 36080 20352 36100
rect 20352 36080 20404 36100
rect 20404 36080 20406 36100
rect 20718 37304 20774 37360
rect 20718 36488 20774 36544
rect 20626 36080 20682 36136
rect 20350 32680 20406 32736
rect 20166 30252 20222 30288
rect 20166 30232 20168 30252
rect 20168 30232 20220 30252
rect 20220 30232 20222 30252
rect 20810 32444 20812 32464
rect 20812 32444 20864 32464
rect 20864 32444 20866 32464
rect 20810 32408 20866 32444
rect 20718 32000 20774 32056
rect 19798 22072 19854 22128
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19890 18828 19946 18864
rect 19890 18808 19892 18828
rect 19892 18808 19944 18828
rect 19944 18808 19946 18828
rect 19890 15564 19946 15600
rect 19890 15544 19892 15564
rect 19892 15544 19944 15564
rect 19944 15544 19946 15564
rect 21270 44820 21272 44840
rect 21272 44820 21324 44840
rect 21324 44820 21326 44840
rect 21270 44784 21326 44820
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22190 52536 22246 52592
rect 21454 35672 21510 35728
rect 21362 32020 21418 32056
rect 21362 32000 21364 32020
rect 21364 32000 21416 32020
rect 21416 32000 21418 32020
rect 21822 41556 21824 41576
rect 21824 41556 21876 41576
rect 21876 41556 21878 41576
rect 21822 41520 21878 41556
rect 21822 37848 21878 37904
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 23202 40976 23258 41032
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 21454 31748 21510 31784
rect 21454 31728 21456 31748
rect 21456 31728 21508 31748
rect 21508 31728 21510 31748
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22190 32428 22246 32464
rect 22190 32408 22192 32428
rect 22192 32408 22244 32428
rect 22244 32408 22246 32428
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22374 32000 22430 32056
rect 22466 31728 22522 31784
rect 22098 26016 22154 26072
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 23754 37576 23810 37632
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22926 31864 22982 31920
rect 23018 31728 23074 31784
rect 22282 25336 22338 25392
rect 22190 19216 22246 19272
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 24030 40296 24086 40352
rect 25134 51856 25190 51912
rect 25042 51176 25098 51232
rect 25042 50496 25098 50552
rect 25042 49816 25098 49872
rect 25042 49172 25044 49192
rect 25044 49172 25096 49192
rect 25096 49172 25098 49192
rect 25042 49136 25098 49172
rect 25042 48456 25098 48512
rect 25042 47776 25098 47832
rect 25042 47096 25098 47152
rect 24766 45736 24822 45792
rect 24674 45056 24730 45112
rect 24858 44396 24914 44432
rect 24858 44376 24860 44396
rect 24860 44376 24912 44396
rect 24912 44376 24914 44396
rect 24858 43016 24914 43072
rect 24766 42336 24822 42392
rect 25318 43696 25374 43752
rect 23938 35672 23994 35728
rect 24858 39616 24914 39672
rect 24858 36896 24914 36952
rect 25134 38936 25190 38992
rect 25318 41656 25374 41712
rect 25318 38256 25374 38312
rect 25410 36216 25466 36272
rect 25318 35536 25374 35592
rect 24030 31456 24086 31512
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 23478 26696 23534 26752
rect 22926 26016 22982 26072
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23386 23296 23442 23352
rect 24122 28736 24178 28792
rect 24398 30504 24454 30560
rect 24490 30368 24546 30424
rect 24858 32852 24860 32872
rect 24860 32852 24912 32872
rect 24912 32852 24914 32872
rect 24858 32816 24914 32852
rect 25502 34856 25558 34912
rect 25410 34176 25466 34232
rect 25318 33496 25374 33552
rect 25134 32716 25136 32736
rect 25136 32716 25188 32736
rect 25188 32716 25190 32736
rect 25134 32680 25190 32716
rect 25318 32136 25374 32192
rect 24858 28056 24914 28112
rect 24950 27376 25006 27432
rect 24766 26016 24822 26072
rect 24950 23976 25006 24032
rect 24950 21956 25006 21992
rect 24950 21936 24952 21956
rect 24952 21936 25004 21956
rect 25004 21936 25006 21956
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17856 23442 17912
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22374 4256 22430 4312
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 24674 21256 24730 21312
rect 24950 20576 25006 20632
rect 24858 19896 24914 19952
rect 25410 30776 25466 30832
rect 25318 30096 25374 30152
rect 25318 29416 25374 29472
rect 25134 24656 25190 24712
rect 26054 22616 26110 22672
rect 23846 18536 23902 18592
rect 23846 17176 23902 17232
rect 24766 16496 24822 16552
rect 24858 15816 24914 15872
rect 25134 15136 25190 15192
rect 24858 14456 24914 14512
rect 24766 13776 24822 13832
rect 24674 13096 24730 13152
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24858 12416 24914 12472
rect 25318 11736 25374 11792
rect 24766 11056 24822 11112
rect 24766 10376 24822 10432
rect 24950 9696 25006 9752
rect 25134 9016 25190 9072
rect 24766 8336 24822 8392
rect 24490 6724 24546 6760
rect 24490 6704 24492 6724
rect 24492 6704 24544 6724
rect 24544 6704 24546 6724
rect 24490 5636 24546 5672
rect 24490 5616 24492 5636
rect 24492 5616 24544 5636
rect 24544 5616 24546 5636
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24766 6976 24822 7032
rect 24950 7656 25006 7712
rect 24950 6296 25006 6352
rect 24766 5616 24822 5672
rect 25318 4936 25374 4992
<< metal3 >>
rect 0 55042 800 55072
rect 2773 55042 2839 55045
rect 0 55040 2839 55042
rect 0 54984 2778 55040
rect 2834 54984 2839 55040
rect 0 54982 2839 54984
rect 0 54952 800 54982
rect 2773 54979 2839 54982
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 14825 53954 14891 53957
rect 14958 53954 14964 53956
rect 14825 53952 14964 53954
rect 14825 53896 14830 53952
rect 14886 53896 14964 53952
rect 14825 53894 14964 53896
rect 14825 53891 14891 53894
rect 14958 53892 14964 53894
rect 15028 53892 15034 53956
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 2946 52800 3262 52801
rect 0 52730 800 52760
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 1301 52730 1367 52733
rect 0 52728 1367 52730
rect 0 52672 1306 52728
rect 1362 52672 1367 52728
rect 0 52670 1367 52672
rect 0 52640 800 52670
rect 1301 52667 1367 52670
rect 14549 52596 14615 52597
rect 14549 52592 14596 52596
rect 14660 52594 14666 52596
rect 22185 52594 22251 52597
rect 22318 52594 22324 52596
rect 14549 52536 14554 52592
rect 14549 52532 14596 52536
rect 14660 52534 14706 52594
rect 22185 52592 22324 52594
rect 22185 52536 22190 52592
rect 22246 52536 22324 52592
rect 22185 52534 22324 52536
rect 14660 52532 14666 52534
rect 14549 52531 14615 52532
rect 22185 52531 22251 52534
rect 22318 52532 22324 52534
rect 22388 52532 22394 52596
rect 26200 52504 27000 52624
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 25129 51914 25195 51917
rect 26200 51914 27000 51944
rect 25129 51912 27000 51914
rect 25129 51856 25134 51912
rect 25190 51856 27000 51912
rect 25129 51854 27000 51856
rect 25129 51851 25195 51854
rect 26200 51824 27000 51854
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25037 51234 25103 51237
rect 26200 51234 27000 51264
rect 25037 51232 27000 51234
rect 25037 51176 25042 51232
rect 25098 51176 27000 51232
rect 25037 51174 27000 51176
rect 25037 51171 25103 51174
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 26200 51144 27000 51174
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 25037 50552 27000 50554
rect 25037 50496 25042 50552
rect 25098 50496 27000 50552
rect 25037 50494 27000 50496
rect 25037 50491 25103 50494
rect 26200 50464 27000 50494
rect 0 50418 800 50448
rect 933 50418 999 50421
rect 0 50416 999 50418
rect 0 50360 938 50416
rect 994 50360 999 50416
rect 0 50358 999 50360
rect 0 50328 800 50358
rect 933 50355 999 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25037 49874 25103 49877
rect 26200 49874 27000 49904
rect 25037 49872 27000 49874
rect 25037 49816 25042 49872
rect 25098 49816 27000 49872
rect 25037 49814 27000 49816
rect 25037 49811 25103 49814
rect 26200 49784 27000 49814
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 25037 49194 25103 49197
rect 26200 49194 27000 49224
rect 25037 49192 27000 49194
rect 25037 49136 25042 49192
rect 25098 49136 27000 49192
rect 25037 49134 27000 49136
rect 25037 49131 25103 49134
rect 26200 49104 27000 49134
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25037 48514 25103 48517
rect 26200 48514 27000 48544
rect 25037 48512 27000 48514
rect 25037 48456 25042 48512
rect 25098 48456 27000 48512
rect 25037 48454 27000 48456
rect 25037 48451 25103 48454
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 26200 48424 27000 48454
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 933 48106 999 48109
rect 0 48104 999 48106
rect 0 48048 938 48104
rect 994 48048 999 48104
rect 0 48046 999 48048
rect 0 48016 800 48046
rect 933 48043 999 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 25037 47834 25103 47837
rect 26200 47834 27000 47864
rect 25037 47832 27000 47834
rect 25037 47776 25042 47832
rect 25098 47776 27000 47832
rect 25037 47774 27000 47776
rect 25037 47771 25103 47774
rect 26200 47744 27000 47774
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25037 47154 25103 47157
rect 26200 47154 27000 47184
rect 25037 47152 27000 47154
rect 25037 47096 25042 47152
rect 25098 47096 27000 47152
rect 25037 47094 27000 47096
rect 25037 47091 25103 47094
rect 26200 47064 27000 47094
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 17166 46412 17172 46476
rect 17236 46474 17242 46476
rect 18413 46474 18479 46477
rect 17236 46472 18479 46474
rect 17236 46416 18418 46472
rect 18474 46416 18479 46472
rect 17236 46414 18479 46416
rect 17236 46412 17242 46414
rect 18413 46411 18479 46414
rect 26200 46384 27000 46504
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 15326 46004 15332 46068
rect 15396 46066 15402 46068
rect 15561 46066 15627 46069
rect 15396 46064 15627 46066
rect 15396 46008 15566 46064
rect 15622 46008 15627 46064
rect 15396 46006 15627 46008
rect 15396 46004 15402 46006
rect 15561 46003 15627 46006
rect 0 45794 800 45824
rect 933 45794 999 45797
rect 19793 45796 19859 45797
rect 0 45792 999 45794
rect 0 45736 938 45792
rect 994 45736 999 45792
rect 0 45734 999 45736
rect 0 45704 800 45734
rect 933 45731 999 45734
rect 19742 45732 19748 45796
rect 19812 45794 19859 45796
rect 24761 45794 24827 45797
rect 26200 45794 27000 45824
rect 19812 45792 19904 45794
rect 19854 45736 19904 45792
rect 19812 45734 19904 45736
rect 24761 45792 27000 45794
rect 24761 45736 24766 45792
rect 24822 45736 27000 45792
rect 24761 45734 27000 45736
rect 19812 45732 19859 45734
rect 19793 45731 19859 45732
rect 24761 45731 24827 45734
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 26200 45704 27000 45734
rect 17946 45663 18262 45664
rect 19374 45596 19380 45660
rect 19444 45658 19450 45660
rect 20621 45658 20687 45661
rect 19444 45656 20687 45658
rect 19444 45600 20626 45656
rect 20682 45600 20687 45656
rect 19444 45598 20687 45600
rect 19444 45596 19450 45598
rect 20621 45595 20687 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 24669 45114 24735 45117
rect 26200 45114 27000 45144
rect 24669 45112 27000 45114
rect 24669 45056 24674 45112
rect 24730 45056 27000 45112
rect 24669 45054 27000 45056
rect 24669 45051 24735 45054
rect 26200 45024 27000 45054
rect 20662 44780 20668 44844
rect 20732 44842 20738 44844
rect 21265 44842 21331 44845
rect 20732 44840 21331 44842
rect 20732 44784 21270 44840
rect 21326 44784 21331 44840
rect 20732 44782 21331 44784
rect 20732 44780 20738 44782
rect 21265 44779 21331 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 24853 44434 24919 44437
rect 26200 44434 27000 44464
rect 24853 44432 27000 44434
rect 24853 44376 24858 44432
rect 24914 44376 27000 44432
rect 24853 44374 27000 44376
rect 24853 44371 24919 44374
rect 26200 44344 27000 44374
rect 7189 44298 7255 44301
rect 11789 44300 11855 44301
rect 10910 44298 10916 44300
rect 7189 44296 10916 44298
rect 7189 44240 7194 44296
rect 7250 44240 10916 44296
rect 7189 44238 10916 44240
rect 7189 44235 7255 44238
rect 10910 44236 10916 44238
rect 10980 44236 10986 44300
rect 11789 44296 11836 44300
rect 11900 44298 11906 44300
rect 11789 44240 11794 44296
rect 11789 44236 11836 44240
rect 11900 44238 11946 44298
rect 11900 44236 11906 44238
rect 11789 44235 11855 44236
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 25313 43754 25379 43757
rect 26200 43754 27000 43784
rect 25313 43752 27000 43754
rect 25313 43696 25318 43752
rect 25374 43696 27000 43752
rect 25313 43694 27000 43696
rect 25313 43691 25379 43694
rect 26200 43664 27000 43694
rect 7946 43552 8262 43553
rect 0 43392 800 43512
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 24853 43074 24919 43077
rect 26200 43074 27000 43104
rect 24853 43072 27000 43074
rect 24853 43016 24858 43072
rect 24914 43016 27000 43072
rect 24853 43014 27000 43016
rect 24853 43011 24919 43014
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 26200 42984 27000 43014
rect 22946 42943 23262 42944
rect 10225 42938 10291 42941
rect 12566 42938 12572 42940
rect 10225 42936 12572 42938
rect 10225 42880 10230 42936
rect 10286 42880 12572 42936
rect 10225 42878 12572 42880
rect 10225 42875 10291 42878
rect 12566 42876 12572 42878
rect 12636 42876 12642 42940
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 24761 42394 24827 42397
rect 26200 42394 27000 42424
rect 24761 42392 27000 42394
rect 24761 42336 24766 42392
rect 24822 42336 27000 42392
rect 24761 42334 27000 42336
rect 24761 42331 24827 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25313 41714 25379 41717
rect 26200 41714 27000 41744
rect 25313 41712 27000 41714
rect 25313 41656 25318 41712
rect 25374 41656 27000 41712
rect 25313 41654 27000 41656
rect 25313 41651 25379 41654
rect 26200 41624 27000 41654
rect 21817 41578 21883 41581
rect 21950 41578 21956 41580
rect 21817 41576 21956 41578
rect 21817 41520 21822 41576
rect 21878 41520 21956 41576
rect 21817 41518 21956 41520
rect 21817 41515 21883 41518
rect 21950 41516 21956 41518
rect 22020 41516 22026 41580
rect 10317 41442 10383 41445
rect 13670 41442 13676 41444
rect 10317 41440 13676 41442
rect 10317 41384 10322 41440
rect 10378 41384 13676 41440
rect 10317 41382 13676 41384
rect 10317 41379 10383 41382
rect 13670 41380 13676 41382
rect 13740 41380 13746 41444
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 0 41170 800 41200
rect 1669 41170 1735 41173
rect 0 41168 1735 41170
rect 0 41112 1674 41168
rect 1730 41112 1735 41168
rect 0 41110 1735 41112
rect 0 41080 800 41110
rect 1669 41107 1735 41110
rect 23197 41034 23263 41037
rect 26200 41034 27000 41064
rect 23197 41032 27000 41034
rect 23197 40976 23202 41032
rect 23258 40976 27000 41032
rect 23197 40974 27000 40976
rect 23197 40971 23263 40974
rect 26200 40944 27000 40974
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 24025 40354 24091 40357
rect 26200 40354 27000 40384
rect 24025 40352 27000 40354
rect 24025 40296 24030 40352
rect 24086 40296 27000 40352
rect 24025 40294 27000 40296
rect 24025 40291 24091 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 26200 40264 27000 40294
rect 17946 40223 18262 40224
rect 17718 40020 17724 40084
rect 17788 40082 17794 40084
rect 19149 40082 19215 40085
rect 17788 40080 19215 40082
rect 17788 40024 19154 40080
rect 19210 40024 19215 40080
rect 17788 40022 19215 40024
rect 17788 40020 17794 40022
rect 19149 40019 19215 40022
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 24853 39674 24919 39677
rect 26200 39674 27000 39704
rect 24853 39672 27000 39674
rect 24853 39616 24858 39672
rect 24914 39616 27000 39672
rect 24853 39614 27000 39616
rect 24853 39611 24919 39614
rect 26200 39584 27000 39614
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25129 38994 25195 38997
rect 26200 38994 27000 39024
rect 25129 38992 27000 38994
rect 25129 38936 25134 38992
rect 25190 38936 27000 38992
rect 25129 38934 27000 38936
rect 25129 38931 25195 38934
rect 26200 38904 27000 38934
rect 0 38858 800 38888
rect 933 38858 999 38861
rect 0 38856 999 38858
rect 0 38800 938 38856
rect 994 38800 999 38856
rect 0 38798 999 38800
rect 0 38768 800 38798
rect 933 38795 999 38798
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 10910 38524 10916 38588
rect 10980 38586 10986 38588
rect 12750 38586 12756 38588
rect 10980 38526 12756 38586
rect 10980 38524 10986 38526
rect 12750 38524 12756 38526
rect 12820 38524 12826 38588
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 13670 38116 13676 38180
rect 13740 38178 13746 38180
rect 16205 38178 16271 38181
rect 13740 38176 16271 38178
rect 13740 38120 16210 38176
rect 16266 38120 16271 38176
rect 13740 38118 16271 38120
rect 13740 38116 13746 38118
rect 16205 38115 16271 38118
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 21817 37906 21883 37909
rect 16806 37904 21883 37906
rect 16806 37848 21822 37904
rect 21878 37848 21883 37904
rect 16806 37846 21883 37848
rect 15142 37708 15148 37772
rect 15212 37770 15218 37772
rect 15285 37770 15351 37773
rect 16806 37770 16866 37846
rect 21817 37843 21883 37846
rect 15212 37768 16866 37770
rect 15212 37712 15290 37768
rect 15346 37712 16866 37768
rect 15212 37710 16866 37712
rect 16941 37770 17007 37773
rect 17350 37770 17356 37772
rect 16941 37768 17356 37770
rect 16941 37712 16946 37768
rect 17002 37712 17356 37768
rect 16941 37710 17356 37712
rect 15212 37708 15218 37710
rect 15285 37707 15351 37710
rect 16941 37707 17007 37710
rect 17350 37708 17356 37710
rect 17420 37770 17426 37772
rect 17861 37770 17927 37773
rect 17420 37768 17927 37770
rect 17420 37712 17866 37768
rect 17922 37712 17927 37768
rect 17420 37710 17927 37712
rect 17420 37708 17426 37710
rect 17861 37707 17927 37710
rect 23749 37634 23815 37637
rect 26200 37634 27000 37664
rect 23749 37632 27000 37634
rect 23749 37576 23754 37632
rect 23810 37576 27000 37632
rect 23749 37574 27000 37576
rect 23749 37571 23815 37574
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 26200 37544 27000 37574
rect 22946 37503 23262 37504
rect 20110 37300 20116 37364
rect 20180 37362 20186 37364
rect 20713 37362 20779 37365
rect 20180 37360 20779 37362
rect 20180 37304 20718 37360
rect 20774 37304 20779 37360
rect 20180 37302 20779 37304
rect 20180 37300 20186 37302
rect 20713 37299 20779 37302
rect 12566 37028 12572 37092
rect 12636 37090 12642 37092
rect 17585 37090 17651 37093
rect 12636 37088 17651 37090
rect 12636 37032 17590 37088
rect 17646 37032 17651 37088
rect 12636 37030 17651 37032
rect 12636 37028 12642 37030
rect 17585 37027 17651 37030
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 24853 36954 24919 36957
rect 26200 36954 27000 36984
rect 24853 36952 27000 36954
rect 24853 36896 24858 36952
rect 24914 36896 27000 36952
rect 24853 36894 27000 36896
rect 24853 36891 24919 36894
rect 26200 36864 27000 36894
rect 16205 36682 16271 36685
rect 18321 36682 18387 36685
rect 16205 36680 18387 36682
rect 16205 36624 16210 36680
rect 16266 36624 18326 36680
rect 18382 36624 18387 36680
rect 16205 36622 18387 36624
rect 16205 36619 16271 36622
rect 18321 36619 18387 36622
rect 18505 36682 18571 36685
rect 18638 36682 18644 36684
rect 18505 36680 18644 36682
rect 18505 36624 18510 36680
rect 18566 36624 18644 36680
rect 18505 36622 18644 36624
rect 18505 36619 18571 36622
rect 18638 36620 18644 36622
rect 18708 36682 18714 36684
rect 18873 36682 18939 36685
rect 18708 36680 18939 36682
rect 18708 36624 18878 36680
rect 18934 36624 18939 36680
rect 18708 36622 18939 36624
rect 18708 36620 18714 36622
rect 18873 36619 18939 36622
rect 0 36546 800 36576
rect 933 36546 999 36549
rect 0 36544 999 36546
rect 0 36488 938 36544
rect 994 36488 999 36544
rect 0 36486 999 36488
rect 0 36456 800 36486
rect 933 36483 999 36486
rect 17585 36546 17651 36549
rect 20713 36546 20779 36549
rect 17585 36544 20779 36546
rect 17585 36488 17590 36544
rect 17646 36488 20718 36544
rect 20774 36488 20779 36544
rect 17585 36486 20779 36488
rect 17585 36483 17651 36486
rect 20713 36483 20779 36486
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 17677 36410 17743 36413
rect 14966 36408 17743 36410
rect 14966 36352 17682 36408
rect 17738 36352 17743 36408
rect 14966 36350 17743 36352
rect 9029 36138 9095 36141
rect 14966 36138 15026 36350
rect 17677 36347 17743 36350
rect 15285 36274 15351 36277
rect 20437 36274 20503 36277
rect 25405 36274 25471 36277
rect 26200 36274 27000 36304
rect 15285 36272 20546 36274
rect 15285 36216 15290 36272
rect 15346 36216 20442 36272
rect 20498 36216 20546 36272
rect 15285 36214 20546 36216
rect 15285 36211 15351 36214
rect 20437 36211 20546 36214
rect 25405 36272 27000 36274
rect 25405 36216 25410 36272
rect 25466 36216 27000 36272
rect 25405 36214 27000 36216
rect 25405 36211 25471 36214
rect 20345 36138 20411 36141
rect 9029 36136 15026 36138
rect 9029 36080 9034 36136
rect 9090 36080 15026 36136
rect 9029 36078 15026 36080
rect 17726 36136 20411 36138
rect 17726 36080 20350 36136
rect 20406 36080 20411 36136
rect 17726 36078 20411 36080
rect 20486 36138 20546 36211
rect 26200 36184 27000 36214
rect 20621 36138 20687 36141
rect 20486 36136 20687 36138
rect 20486 36080 20626 36136
rect 20682 36080 20687 36136
rect 20486 36078 20687 36080
rect 9029 36075 9095 36078
rect 11881 36004 11947 36005
rect 11830 36002 11836 36004
rect 11790 35942 11836 36002
rect 11900 36002 11947 36004
rect 17726 36002 17786 36078
rect 20345 36075 20411 36078
rect 20621 36075 20687 36078
rect 11900 36000 17786 36002
rect 11942 35944 17786 36000
rect 11830 35940 11836 35942
rect 11900 35942 17786 35944
rect 11900 35940 11947 35942
rect 11881 35939 11947 35940
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 18597 35730 18663 35733
rect 21449 35730 21515 35733
rect 23933 35730 23999 35733
rect 18597 35728 23999 35730
rect 18597 35672 18602 35728
rect 18658 35672 21454 35728
rect 21510 35672 23938 35728
rect 23994 35672 23999 35728
rect 18597 35670 23999 35672
rect 18597 35667 18663 35670
rect 21449 35667 21515 35670
rect 23933 35667 23999 35670
rect 25313 35594 25379 35597
rect 26200 35594 27000 35624
rect 25313 35592 27000 35594
rect 25313 35536 25318 35592
rect 25374 35536 27000 35592
rect 25313 35534 27000 35536
rect 25313 35531 25379 35534
rect 26200 35504 27000 35534
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 12750 35124 12756 35188
rect 12820 35186 12826 35188
rect 13629 35186 13695 35189
rect 12820 35184 13695 35186
rect 12820 35128 13634 35184
rect 13690 35128 13695 35184
rect 12820 35126 13695 35128
rect 12820 35124 12826 35126
rect 13629 35123 13695 35126
rect 25497 34914 25563 34917
rect 26200 34914 27000 34944
rect 25497 34912 27000 34914
rect 25497 34856 25502 34912
rect 25558 34856 27000 34912
rect 25497 34854 27000 34856
rect 25497 34851 25563 34854
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 26200 34824 27000 34854
rect 17946 34783 18262 34784
rect 10869 34642 10935 34645
rect 19517 34642 19583 34645
rect 10869 34640 19583 34642
rect 10869 34584 10874 34640
rect 10930 34584 19522 34640
rect 19578 34584 19583 34640
rect 10869 34582 19583 34584
rect 10869 34579 10935 34582
rect 19517 34579 19583 34582
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 1761 34234 1827 34237
rect 0 34232 1827 34234
rect 0 34176 1766 34232
rect 1822 34176 1827 34232
rect 0 34174 1827 34176
rect 0 34144 800 34174
rect 1761 34171 1827 34174
rect 25405 34234 25471 34237
rect 26200 34234 27000 34264
rect 25405 34232 27000 34234
rect 25405 34176 25410 34232
rect 25466 34176 27000 34232
rect 25405 34174 27000 34176
rect 25405 34171 25471 34174
rect 26200 34144 27000 34174
rect 11881 33826 11947 33829
rect 12198 33826 12204 33828
rect 11881 33824 12204 33826
rect 11881 33768 11886 33824
rect 11942 33768 12204 33824
rect 11881 33766 12204 33768
rect 11881 33763 11947 33766
rect 12198 33764 12204 33766
rect 12268 33764 12274 33828
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33554 25379 33557
rect 26200 33554 27000 33584
rect 25313 33552 27000 33554
rect 25313 33496 25318 33552
rect 25374 33496 27000 33552
rect 25313 33494 27000 33496
rect 25313 33491 25379 33494
rect 26200 33464 27000 33494
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 24853 32874 24919 32877
rect 26200 32874 27000 32904
rect 24853 32872 27000 32874
rect 24853 32816 24858 32872
rect 24914 32816 27000 32872
rect 24853 32814 27000 32816
rect 24853 32811 24919 32814
rect 26200 32784 27000 32814
rect 20345 32738 20411 32741
rect 25129 32738 25195 32741
rect 20345 32736 25195 32738
rect 20345 32680 20350 32736
rect 20406 32680 25134 32736
rect 25190 32680 25195 32736
rect 20345 32678 25195 32680
rect 20345 32675 20411 32678
rect 25129 32675 25195 32678
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 17166 32540 17172 32604
rect 17236 32602 17242 32604
rect 17309 32602 17375 32605
rect 17236 32600 17375 32602
rect 17236 32544 17314 32600
rect 17370 32544 17375 32600
rect 17236 32542 17375 32544
rect 17236 32540 17242 32542
rect 17309 32539 17375 32542
rect 14590 32404 14596 32468
rect 14660 32466 14666 32468
rect 16757 32466 16823 32469
rect 14660 32464 16823 32466
rect 14660 32408 16762 32464
rect 16818 32408 16823 32464
rect 14660 32406 16823 32408
rect 14660 32404 14666 32406
rect 16757 32403 16823 32406
rect 20805 32466 20871 32469
rect 22185 32466 22251 32469
rect 20805 32464 22251 32466
rect 20805 32408 20810 32464
rect 20866 32408 22190 32464
rect 22246 32408 22251 32464
rect 20805 32406 22251 32408
rect 20805 32403 20871 32406
rect 22185 32403 22251 32406
rect 17033 32194 17099 32197
rect 17677 32194 17743 32197
rect 17033 32192 17743 32194
rect 17033 32136 17038 32192
rect 17094 32136 17682 32192
rect 17738 32136 17743 32192
rect 17033 32134 17743 32136
rect 17033 32131 17099 32134
rect 17677 32131 17743 32134
rect 25313 32194 25379 32197
rect 26200 32194 27000 32224
rect 25313 32192 27000 32194
rect 25313 32136 25318 32192
rect 25374 32136 27000 32192
rect 25313 32134 27000 32136
rect 25313 32131 25379 32134
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 26200 32104 27000 32134
rect 22946 32063 23262 32064
rect 14273 32058 14339 32061
rect 20110 32058 20116 32060
rect 14273 32056 20116 32058
rect 14273 32000 14278 32056
rect 14334 32000 20116 32056
rect 14273 31998 20116 32000
rect 14273 31995 14339 31998
rect 20110 31996 20116 31998
rect 20180 31996 20186 32060
rect 20713 32058 20779 32061
rect 21357 32058 21423 32061
rect 20713 32056 21423 32058
rect 20713 32000 20718 32056
rect 20774 32000 21362 32056
rect 21418 32000 21423 32056
rect 20713 31998 21423 32000
rect 20713 31995 20779 31998
rect 21357 31995 21423 31998
rect 22369 32058 22435 32061
rect 22369 32056 22570 32058
rect 22369 32000 22374 32056
rect 22430 32000 22570 32056
rect 22369 31998 22570 32000
rect 22369 31995 22435 31998
rect 0 31922 800 31952
rect 933 31922 999 31925
rect 0 31920 999 31922
rect 0 31864 938 31920
rect 994 31864 999 31920
rect 0 31862 999 31864
rect 0 31832 800 31862
rect 933 31859 999 31862
rect 9029 31922 9095 31925
rect 9397 31922 9463 31925
rect 9029 31920 9463 31922
rect 9029 31864 9034 31920
rect 9090 31864 9402 31920
rect 9458 31864 9463 31920
rect 9029 31862 9463 31864
rect 22510 31922 22570 31998
rect 22921 31922 22987 31925
rect 22510 31920 22987 31922
rect 22510 31864 22926 31920
rect 22982 31864 22987 31920
rect 22510 31862 22987 31864
rect 9029 31859 9095 31862
rect 9397 31859 9463 31862
rect 22921 31859 22987 31862
rect 15142 31724 15148 31788
rect 15212 31786 15218 31788
rect 19926 31786 19932 31788
rect 15212 31726 19932 31786
rect 15212 31724 15218 31726
rect 19926 31724 19932 31726
rect 19996 31724 20002 31788
rect 21449 31786 21515 31789
rect 22318 31786 22324 31788
rect 21449 31784 22324 31786
rect 21449 31728 21454 31784
rect 21510 31728 22324 31784
rect 21449 31726 22324 31728
rect 21449 31723 21515 31726
rect 22318 31724 22324 31726
rect 22388 31724 22394 31788
rect 22461 31786 22527 31789
rect 23013 31786 23079 31789
rect 22461 31784 23079 31786
rect 22461 31728 22466 31784
rect 22522 31728 23018 31784
rect 23074 31728 23079 31784
rect 22461 31726 23079 31728
rect 22461 31723 22527 31726
rect 23013 31723 23079 31726
rect 12709 31650 12775 31653
rect 13670 31650 13676 31652
rect 12709 31648 13676 31650
rect 12709 31592 12714 31648
rect 12770 31592 13676 31648
rect 12709 31590 13676 31592
rect 12709 31587 12775 31590
rect 13670 31588 13676 31590
rect 13740 31588 13746 31652
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 24025 31514 24091 31517
rect 26200 31514 27000 31544
rect 24025 31512 27000 31514
rect 24025 31456 24030 31512
rect 24086 31456 27000 31512
rect 24025 31454 27000 31456
rect 24025 31451 24091 31454
rect 26200 31424 27000 31454
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25405 30834 25471 30837
rect 26200 30834 27000 30864
rect 25405 30832 27000 30834
rect 25405 30776 25410 30832
rect 25466 30776 27000 30832
rect 25405 30774 27000 30776
rect 25405 30771 25471 30774
rect 26200 30744 27000 30774
rect 13353 30562 13419 30565
rect 24393 30564 24459 30565
rect 13486 30562 13492 30564
rect 13353 30560 13492 30562
rect 13353 30504 13358 30560
rect 13414 30504 13492 30560
rect 13353 30502 13492 30504
rect 13353 30499 13419 30502
rect 13486 30500 13492 30502
rect 13556 30500 13562 30564
rect 24342 30562 24348 30564
rect 24302 30502 24348 30562
rect 24412 30560 24459 30564
rect 24454 30504 24459 30560
rect 24342 30500 24348 30502
rect 24412 30500 24459 30504
rect 24393 30499 24459 30500
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 24485 30428 24551 30429
rect 24485 30424 24532 30428
rect 24596 30426 24602 30428
rect 24485 30368 24490 30424
rect 24485 30364 24532 30368
rect 24596 30366 24642 30426
rect 24596 30364 24602 30366
rect 24485 30363 24551 30364
rect 19149 30290 19215 30293
rect 19374 30290 19380 30292
rect 19149 30288 19380 30290
rect 19149 30232 19154 30288
rect 19210 30232 19380 30288
rect 19149 30230 19380 30232
rect 19149 30227 19215 30230
rect 19374 30228 19380 30230
rect 19444 30228 19450 30292
rect 19742 30228 19748 30292
rect 19812 30290 19818 30292
rect 20161 30290 20227 30293
rect 19812 30288 20227 30290
rect 19812 30232 20166 30288
rect 20222 30232 20227 30288
rect 19812 30230 20227 30232
rect 19812 30228 19818 30230
rect 20161 30227 20227 30230
rect 12566 30092 12572 30156
rect 12636 30154 12642 30156
rect 12985 30154 13051 30157
rect 12636 30152 13051 30154
rect 12636 30096 12990 30152
rect 13046 30096 13051 30152
rect 12636 30094 13051 30096
rect 12636 30092 12642 30094
rect 12985 30091 13051 30094
rect 15285 30154 15351 30157
rect 15510 30154 15516 30156
rect 15285 30152 15516 30154
rect 15285 30096 15290 30152
rect 15346 30096 15516 30152
rect 15285 30094 15516 30096
rect 15285 30091 15351 30094
rect 15510 30092 15516 30094
rect 15580 30092 15586 30156
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 0 29610 800 29640
rect 1301 29610 1367 29613
rect 0 29608 1367 29610
rect 0 29552 1306 29608
rect 1362 29552 1367 29608
rect 0 29550 1367 29552
rect 0 29520 800 29550
rect 1301 29547 1367 29550
rect 17585 29476 17651 29477
rect 17534 29412 17540 29476
rect 17604 29474 17651 29476
rect 25313 29474 25379 29477
rect 26200 29474 27000 29504
rect 17604 29472 17696 29474
rect 17646 29416 17696 29472
rect 17604 29414 17696 29416
rect 25313 29472 27000 29474
rect 25313 29416 25318 29472
rect 25374 29416 27000 29472
rect 25313 29414 27000 29416
rect 17604 29412 17651 29414
rect 17585 29411 17651 29412
rect 25313 29411 25379 29414
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 26200 29384 27000 29414
rect 17946 29343 18262 29344
rect 18965 29338 19031 29341
rect 19517 29338 19583 29341
rect 18965 29336 19583 29338
rect 18965 29280 18970 29336
rect 19026 29280 19522 29336
rect 19578 29280 19583 29336
rect 18965 29278 19583 29280
rect 18965 29275 19031 29278
rect 19517 29275 19583 29278
rect 15510 29004 15516 29068
rect 15580 29066 15586 29068
rect 16481 29066 16547 29069
rect 15580 29064 16547 29066
rect 15580 29008 16486 29064
rect 16542 29008 16547 29064
rect 15580 29006 16547 29008
rect 15580 29004 15586 29006
rect 16481 29003 16547 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24117 28794 24183 28797
rect 26200 28794 27000 28824
rect 24117 28792 27000 28794
rect 24117 28736 24122 28792
rect 24178 28736 27000 28792
rect 24117 28734 27000 28736
rect 24117 28731 24183 28734
rect 26200 28704 27000 28734
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 24853 28114 24919 28117
rect 26200 28114 27000 28144
rect 24853 28112 27000 28114
rect 24853 28056 24858 28112
rect 24914 28056 27000 28112
rect 24853 28054 27000 28056
rect 24853 28051 24919 28054
rect 26200 28024 27000 28054
rect 12065 27978 12131 27981
rect 18413 27978 18479 27981
rect 18873 27978 18939 27981
rect 12065 27976 18939 27978
rect 12065 27920 12070 27976
rect 12126 27920 18418 27976
rect 18474 27920 18878 27976
rect 18934 27920 18939 27976
rect 12065 27918 18939 27920
rect 12065 27915 12131 27918
rect 18413 27915 18479 27918
rect 18873 27915 18939 27918
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 14958 27570 14964 27572
rect 12390 27510 14964 27570
rect 12249 27434 12315 27437
rect 12390 27434 12450 27510
rect 14958 27508 14964 27510
rect 15028 27570 15034 27572
rect 17953 27570 18019 27573
rect 18413 27572 18479 27573
rect 18413 27570 18460 27572
rect 15028 27568 18019 27570
rect 15028 27512 17958 27568
rect 18014 27512 18019 27568
rect 15028 27510 18019 27512
rect 18372 27568 18460 27570
rect 18524 27570 18530 27572
rect 21950 27570 21956 27572
rect 18372 27512 18418 27568
rect 18372 27510 18460 27512
rect 15028 27508 15034 27510
rect 17953 27507 18019 27510
rect 18413 27508 18460 27510
rect 18524 27510 21956 27570
rect 18524 27508 18530 27510
rect 21950 27508 21956 27510
rect 22020 27508 22026 27572
rect 18413 27507 18479 27508
rect 12249 27432 12450 27434
rect 12249 27376 12254 27432
rect 12310 27376 12450 27432
rect 12249 27374 12450 27376
rect 17861 27434 17927 27437
rect 20662 27434 20668 27436
rect 17861 27432 20668 27434
rect 17861 27376 17866 27432
rect 17922 27376 20668 27432
rect 17861 27374 20668 27376
rect 12249 27371 12315 27374
rect 17861 27371 17927 27374
rect 20662 27372 20668 27374
rect 20732 27372 20738 27436
rect 24945 27434 25011 27437
rect 26200 27434 27000 27464
rect 24945 27432 27000 27434
rect 24945 27376 24950 27432
rect 25006 27376 27000 27432
rect 24945 27374 27000 27376
rect 24945 27371 25011 27374
rect 26200 27344 27000 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 10041 27298 10107 27301
rect 13169 27298 13235 27301
rect 10041 27296 13235 27298
rect 10041 27240 10046 27296
rect 10102 27240 13174 27296
rect 13230 27240 13235 27296
rect 10041 27238 13235 27240
rect 10041 27235 10107 27238
rect 13169 27235 13235 27238
rect 15326 27236 15332 27300
rect 15396 27298 15402 27300
rect 16021 27298 16087 27301
rect 15396 27296 16087 27298
rect 15396 27240 16026 27296
rect 16082 27240 16087 27296
rect 15396 27238 16087 27240
rect 15396 27236 15402 27238
rect 16021 27235 16087 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 14958 26828 14964 26892
rect 15028 26890 15034 26892
rect 15101 26890 15167 26893
rect 15028 26888 15167 26890
rect 15028 26832 15106 26888
rect 15162 26832 15167 26888
rect 15028 26830 15167 26832
rect 15028 26828 15034 26830
rect 15101 26827 15167 26830
rect 23473 26754 23539 26757
rect 26200 26754 27000 26784
rect 23473 26752 27000 26754
rect 23473 26696 23478 26752
rect 23534 26696 27000 26752
rect 23473 26694 27000 26696
rect 23473 26691 23539 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 26200 26664 27000 26694
rect 22946 26623 23262 26624
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 22093 26074 22159 26077
rect 22921 26074 22987 26077
rect 22093 26072 22987 26074
rect 22093 26016 22098 26072
rect 22154 26016 22926 26072
rect 22982 26016 22987 26072
rect 22093 26014 22987 26016
rect 22093 26011 22159 26014
rect 22921 26011 22987 26014
rect 24761 26074 24827 26077
rect 26200 26074 27000 26104
rect 24761 26072 27000 26074
rect 24761 26016 24766 26072
rect 24822 26016 27000 26072
rect 24761 26014 27000 26016
rect 24761 26011 24827 26014
rect 26200 25984 27000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 22277 25394 22343 25397
rect 26200 25394 27000 25424
rect 22277 25392 27000 25394
rect 22277 25336 22282 25392
rect 22338 25336 27000 25392
rect 22277 25334 27000 25336
rect 22277 25331 22343 25334
rect 26200 25304 27000 25334
rect 12433 25258 12499 25261
rect 12801 25258 12867 25261
rect 12433 25256 12867 25258
rect 12433 25200 12438 25256
rect 12494 25200 12806 25256
rect 12862 25200 12867 25256
rect 12433 25198 12867 25200
rect 12433 25195 12499 25198
rect 12801 25195 12867 25198
rect 12893 25122 12959 25125
rect 14590 25122 14596 25124
rect 12893 25120 14596 25122
rect 12893 25064 12898 25120
rect 12954 25064 14596 25120
rect 12893 25062 14596 25064
rect 12893 25059 12959 25062
rect 14590 25060 14596 25062
rect 14660 25060 14666 25124
rect 7946 25056 8262 25057
rect 0 24986 800 25016
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 1301 24986 1367 24989
rect 0 24984 1367 24986
rect 0 24928 1306 24984
rect 1362 24928 1367 24984
rect 0 24926 1367 24928
rect 0 24896 800 24926
rect 1301 24923 1367 24926
rect 12065 24986 12131 24989
rect 15142 24986 15148 24988
rect 12065 24984 15148 24986
rect 12065 24928 12070 24984
rect 12126 24928 15148 24984
rect 12065 24926 15148 24928
rect 12065 24923 12131 24926
rect 15142 24924 15148 24926
rect 15212 24924 15218 24988
rect 16665 24850 16731 24853
rect 17166 24850 17172 24852
rect 16665 24848 17172 24850
rect 16665 24792 16670 24848
rect 16726 24792 17172 24848
rect 16665 24790 17172 24792
rect 16665 24787 16731 24790
rect 17166 24788 17172 24790
rect 17236 24788 17242 24852
rect 25129 24714 25195 24717
rect 26200 24714 27000 24744
rect 25129 24712 27000 24714
rect 25129 24656 25134 24712
rect 25190 24656 27000 24712
rect 25129 24654 27000 24656
rect 25129 24651 25195 24654
rect 26200 24624 27000 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24945 24034 25011 24037
rect 26200 24034 27000 24064
rect 24945 24032 27000 24034
rect 24945 23976 24950 24032
rect 25006 23976 27000 24032
rect 24945 23974 27000 23976
rect 24945 23971 25011 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 26200 23944 27000 23974
rect 17946 23903 18262 23904
rect 17585 23492 17651 23493
rect 17534 23490 17540 23492
rect 17494 23430 17540 23490
rect 17604 23488 17651 23492
rect 17646 23432 17651 23488
rect 17534 23428 17540 23430
rect 17604 23428 17651 23432
rect 17585 23427 17651 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 23381 23354 23447 23357
rect 26200 23354 27000 23384
rect 23381 23352 27000 23354
rect 23381 23296 23386 23352
rect 23442 23296 27000 23352
rect 23381 23294 27000 23296
rect 23381 23291 23447 23294
rect 26200 23264 27000 23294
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 0 22674 800 22704
rect 1301 22674 1367 22677
rect 0 22672 1367 22674
rect 0 22616 1306 22672
rect 1362 22616 1367 22672
rect 0 22614 1367 22616
rect 0 22584 800 22614
rect 1301 22611 1367 22614
rect 26049 22674 26115 22677
rect 26200 22674 27000 22704
rect 26049 22672 27000 22674
rect 26049 22616 26054 22672
rect 26110 22616 27000 22672
rect 26049 22614 27000 22616
rect 26049 22611 26115 22614
rect 26200 22584 27000 22614
rect 11646 22476 11652 22540
rect 11716 22538 11722 22540
rect 12893 22538 12959 22541
rect 11716 22536 12959 22538
rect 11716 22480 12898 22536
rect 12954 22480 12959 22536
rect 11716 22478 12959 22480
rect 11716 22476 11722 22478
rect 12893 22475 12959 22478
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 16941 22266 17007 22269
rect 17125 22266 17191 22269
rect 16941 22264 17191 22266
rect 16941 22208 16946 22264
rect 17002 22208 17130 22264
rect 17186 22208 17191 22264
rect 16941 22206 17191 22208
rect 16941 22203 17007 22206
rect 17125 22203 17191 22206
rect 17493 22130 17559 22133
rect 19793 22130 19859 22133
rect 17493 22128 19859 22130
rect 17493 22072 17498 22128
rect 17554 22072 19798 22128
rect 19854 22072 19859 22128
rect 17493 22070 19859 22072
rect 17493 22067 17559 22070
rect 19793 22067 19859 22070
rect 12065 21994 12131 21997
rect 17861 21994 17927 21997
rect 12065 21992 17927 21994
rect 12065 21936 12070 21992
rect 12126 21936 17866 21992
rect 17922 21936 17927 21992
rect 12065 21934 17927 21936
rect 12065 21931 12131 21934
rect 17861 21931 17927 21934
rect 24945 21994 25011 21997
rect 26200 21994 27000 22024
rect 24945 21992 27000 21994
rect 24945 21936 24950 21992
rect 25006 21936 27000 21992
rect 24945 21934 27000 21936
rect 24945 21931 25011 21934
rect 26200 21904 27000 21934
rect 12341 21858 12407 21861
rect 15561 21858 15627 21861
rect 12341 21856 15627 21858
rect 12341 21800 12346 21856
rect 12402 21800 15566 21856
rect 15622 21800 15627 21856
rect 12341 21798 15627 21800
rect 12341 21795 12407 21798
rect 15561 21795 15627 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 15510 21660 15516 21724
rect 15580 21722 15586 21724
rect 16113 21722 16179 21725
rect 15580 21720 16179 21722
rect 15580 21664 16118 21720
rect 16174 21664 16179 21720
rect 15580 21662 16179 21664
rect 15580 21660 15586 21662
rect 16113 21659 16179 21662
rect 13486 21524 13492 21588
rect 13556 21586 13562 21588
rect 13905 21586 13971 21589
rect 13556 21584 13971 21586
rect 13556 21528 13910 21584
rect 13966 21528 13971 21584
rect 13556 21526 13971 21528
rect 13556 21524 13562 21526
rect 13905 21523 13971 21526
rect 10409 21450 10475 21453
rect 10542 21450 10548 21452
rect 10409 21448 10548 21450
rect 10409 21392 10414 21448
rect 10470 21392 10548 21448
rect 10409 21390 10548 21392
rect 10409 21387 10475 21390
rect 10542 21388 10548 21390
rect 10612 21388 10618 21452
rect 13445 21450 13511 21453
rect 14549 21450 14615 21453
rect 13445 21448 14615 21450
rect 13445 21392 13450 21448
rect 13506 21392 14554 21448
rect 14610 21392 14615 21448
rect 13445 21390 14615 21392
rect 13445 21387 13511 21390
rect 14549 21387 14615 21390
rect 24669 21314 24735 21317
rect 26200 21314 27000 21344
rect 24669 21312 27000 21314
rect 24669 21256 24674 21312
rect 24730 21256 27000 21312
rect 24669 21254 27000 21256
rect 24669 21251 24735 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 26200 21224 27000 21254
rect 22946 21183 23262 21184
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 17309 20636 17375 20637
rect 17309 20632 17356 20636
rect 17420 20634 17426 20636
rect 24945 20634 25011 20637
rect 26200 20634 27000 20664
rect 17309 20576 17314 20632
rect 17309 20572 17356 20576
rect 17420 20574 17466 20634
rect 24945 20632 27000 20634
rect 24945 20576 24950 20632
rect 25006 20576 27000 20632
rect 24945 20574 27000 20576
rect 17420 20572 17426 20574
rect 17309 20571 17375 20572
rect 24945 20571 25011 20574
rect 26200 20544 27000 20574
rect 17217 20498 17283 20501
rect 18638 20498 18644 20500
rect 17217 20496 18644 20498
rect 17217 20440 17222 20496
rect 17278 20440 18644 20496
rect 17217 20438 18644 20440
rect 17217 20435 17283 20438
rect 18638 20436 18644 20438
rect 18708 20436 18714 20500
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 24853 19954 24919 19957
rect 26200 19954 27000 19984
rect 24853 19952 27000 19954
rect 24853 19896 24858 19952
rect 24914 19896 27000 19952
rect 24853 19894 27000 19896
rect 24853 19891 24919 19894
rect 26200 19864 27000 19894
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 17033 19410 17099 19413
rect 18454 19410 18460 19412
rect 17033 19408 18460 19410
rect 17033 19352 17038 19408
rect 17094 19352 18460 19408
rect 17033 19350 18460 19352
rect 17033 19347 17099 19350
rect 18454 19348 18460 19350
rect 18524 19410 18530 19412
rect 18781 19410 18847 19413
rect 18524 19408 18847 19410
rect 18524 19352 18786 19408
rect 18842 19352 18847 19408
rect 18524 19350 18847 19352
rect 18524 19348 18530 19350
rect 18781 19347 18847 19350
rect 22185 19274 22251 19277
rect 26200 19274 27000 19304
rect 22185 19272 27000 19274
rect 22185 19216 22190 19272
rect 22246 19216 27000 19272
rect 22185 19214 27000 19216
rect 22185 19211 22251 19214
rect 26200 19184 27000 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 19885 18866 19951 18869
rect 20110 18866 20116 18868
rect 19885 18864 20116 18866
rect 19885 18808 19890 18864
rect 19946 18808 20116 18864
rect 19885 18806 20116 18808
rect 19885 18803 19951 18806
rect 20110 18804 20116 18806
rect 20180 18804 20186 18868
rect 23841 18594 23907 18597
rect 26200 18594 27000 18624
rect 23841 18592 27000 18594
rect 23841 18536 23846 18592
rect 23902 18536 27000 18592
rect 23841 18534 27000 18536
rect 23841 18531 23907 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 26200 18504 27000 18534
rect 17946 18463 18262 18464
rect 12198 18396 12204 18460
rect 12268 18458 12274 18460
rect 12341 18458 12407 18461
rect 12268 18456 12407 18458
rect 12268 18400 12346 18456
rect 12402 18400 12407 18456
rect 12268 18398 12407 18400
rect 12268 18396 12274 18398
rect 12341 18395 12407 18398
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 23841 17234 23907 17237
rect 26200 17234 27000 17264
rect 23841 17232 27000 17234
rect 23841 17176 23846 17232
rect 23902 17176 27000 17232
rect 23841 17174 27000 17176
rect 23841 17171 23907 17174
rect 26200 17144 27000 17174
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 15377 16556 15443 16557
rect 15326 16554 15332 16556
rect 15286 16494 15332 16554
rect 15396 16552 15443 16556
rect 15438 16496 15443 16552
rect 15326 16492 15332 16494
rect 15396 16492 15443 16496
rect 15377 16491 15443 16492
rect 24761 16554 24827 16557
rect 26200 16554 27000 16584
rect 24761 16552 27000 16554
rect 24761 16496 24766 16552
rect 24822 16496 27000 16552
rect 24761 16494 27000 16496
rect 24761 16491 24827 16494
rect 26200 16464 27000 16494
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 13997 16282 14063 16285
rect 14958 16282 14964 16284
rect 13997 16280 14964 16282
rect 13997 16224 14002 16280
rect 14058 16224 14964 16280
rect 13997 16222 14964 16224
rect 13997 16219 14063 16222
rect 14958 16220 14964 16222
rect 15028 16282 15034 16284
rect 15193 16282 15259 16285
rect 15028 16280 15259 16282
rect 15028 16224 15198 16280
rect 15254 16224 15259 16280
rect 15028 16222 15259 16224
rect 15028 16220 15034 16222
rect 15193 16219 15259 16222
rect 24853 15874 24919 15877
rect 26200 15874 27000 15904
rect 24853 15872 27000 15874
rect 24853 15816 24858 15872
rect 24914 15816 27000 15872
rect 24853 15814 27000 15816
rect 24853 15811 24919 15814
rect 2946 15808 3262 15809
rect 0 15738 800 15768
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 19885 15604 19951 15605
rect 19885 15602 19932 15604
rect 19840 15600 19932 15602
rect 19840 15544 19890 15600
rect 19840 15542 19932 15544
rect 19885 15540 19932 15542
rect 19996 15540 20002 15604
rect 19885 15539 19951 15540
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 25129 15194 25195 15197
rect 26200 15194 27000 15224
rect 25129 15192 27000 15194
rect 25129 15136 25134 15192
rect 25190 15136 27000 15192
rect 25129 15134 27000 15136
rect 25129 15131 25195 15134
rect 26200 15104 27000 15134
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14514 24919 14517
rect 26200 14514 27000 14544
rect 24853 14512 27000 14514
rect 24853 14456 24858 14512
rect 24914 14456 27000 14512
rect 24853 14454 27000 14456
rect 24853 14451 24919 14454
rect 26200 14424 27000 14454
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 0 13426 800 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 800 13366
rect 2773 13363 2839 13366
rect 24669 13154 24735 13157
rect 26200 13154 27000 13184
rect 24669 13152 27000 13154
rect 24669 13096 24674 13152
rect 24730 13096 27000 13152
rect 24669 13094 27000 13096
rect 24669 13091 24735 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 26200 13064 27000 13094
rect 17946 13023 18262 13024
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 24853 12474 24919 12477
rect 26200 12474 27000 12504
rect 24853 12472 27000 12474
rect 24853 12416 24858 12472
rect 24914 12416 27000 12472
rect 24853 12414 27000 12416
rect 24853 12411 24919 12414
rect 26200 12384 27000 12414
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 25313 11794 25379 11797
rect 26200 11794 27000 11824
rect 25313 11792 27000 11794
rect 25313 11736 25318 11792
rect 25374 11736 27000 11792
rect 25313 11734 27000 11736
rect 25313 11731 25379 11734
rect 26200 11704 27000 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 0 11114 800 11144
rect 2773 11114 2839 11117
rect 0 11112 2839 11114
rect 0 11056 2778 11112
rect 2834 11056 2839 11112
rect 0 11054 2839 11056
rect 0 11024 800 11054
rect 2773 11051 2839 11054
rect 24761 11114 24827 11117
rect 26200 11114 27000 11144
rect 24761 11112 27000 11114
rect 24761 11056 24766 11112
rect 24822 11056 27000 11112
rect 24761 11054 27000 11056
rect 24761 11051 24827 11054
rect 26200 11024 27000 11054
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24761 10434 24827 10437
rect 26200 10434 27000 10464
rect 24761 10432 27000 10434
rect 24761 10376 24766 10432
rect 24822 10376 27000 10432
rect 24761 10374 27000 10376
rect 24761 10371 24827 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 26200 10344 27000 10374
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24945 9754 25011 9757
rect 26200 9754 27000 9784
rect 24945 9752 27000 9754
rect 24945 9696 24950 9752
rect 25006 9696 27000 9752
rect 24945 9694 27000 9696
rect 24945 9691 25011 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 25129 9074 25195 9077
rect 26200 9074 27000 9104
rect 25129 9072 27000 9074
rect 25129 9016 25134 9072
rect 25190 9016 27000 9072
rect 25129 9014 27000 9016
rect 25129 9011 25195 9014
rect 26200 8984 27000 9014
rect 0 8802 800 8832
rect 3049 8802 3115 8805
rect 0 8800 3115 8802
rect 0 8744 3054 8800
rect 3110 8744 3115 8800
rect 0 8742 3115 8744
rect 0 8712 800 8742
rect 3049 8739 3115 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24761 8394 24827 8397
rect 26200 8394 27000 8424
rect 24761 8392 27000 8394
rect 24761 8336 24766 8392
rect 24822 8336 27000 8392
rect 24761 8334 27000 8336
rect 24761 8331 24827 8334
rect 26200 8304 27000 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 7714 25011 7717
rect 26200 7714 27000 7744
rect 24945 7712 27000 7714
rect 24945 7656 24950 7712
rect 25006 7656 27000 7712
rect 24945 7654 27000 7656
rect 24945 7651 25011 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24761 7034 24827 7037
rect 26200 7034 27000 7064
rect 24761 7032 27000 7034
rect 24761 6976 24766 7032
rect 24822 6976 27000 7032
rect 24761 6974 27000 6976
rect 24761 6971 24827 6974
rect 26200 6944 27000 6974
rect 24485 6764 24551 6765
rect 24485 6760 24532 6764
rect 24596 6762 24602 6764
rect 24485 6704 24490 6760
rect 24485 6700 24532 6704
rect 24596 6702 24642 6762
rect 24596 6700 24602 6702
rect 24485 6699 24551 6700
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3141 6490 3207 6493
rect 0 6488 3207 6490
rect 0 6432 3146 6488
rect 3202 6432 3207 6488
rect 0 6430 3207 6432
rect 0 6400 800 6430
rect 3141 6427 3207 6430
rect 24945 6354 25011 6357
rect 26200 6354 27000 6384
rect 24945 6352 27000 6354
rect 24945 6296 24950 6352
rect 25006 6296 27000 6352
rect 24945 6294 27000 6296
rect 24945 6291 25011 6294
rect 26200 6264 27000 6294
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 7833 5674 7899 5677
rect 13486 5674 13492 5676
rect 7833 5672 13492 5674
rect 7833 5616 7838 5672
rect 7894 5616 13492 5672
rect 7833 5614 13492 5616
rect 7833 5611 7899 5614
rect 13486 5612 13492 5614
rect 13556 5612 13562 5676
rect 24342 5612 24348 5676
rect 24412 5674 24418 5676
rect 24485 5674 24551 5677
rect 24412 5672 24551 5674
rect 24412 5616 24490 5672
rect 24546 5616 24551 5672
rect 24412 5614 24551 5616
rect 24412 5612 24418 5614
rect 24485 5611 24551 5614
rect 24761 5674 24827 5677
rect 26200 5674 27000 5704
rect 24761 5672 27000 5674
rect 24761 5616 24766 5672
rect 24822 5616 27000 5672
rect 24761 5614 27000 5616
rect 24761 5611 24827 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 25313 4994 25379 4997
rect 26200 4994 27000 5024
rect 25313 4992 27000 4994
rect 25313 4936 25318 4992
rect 25374 4936 27000 4992
rect 25313 4934 27000 4936
rect 25313 4931 25379 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 26200 4904 27000 4934
rect 22946 4863 23262 4864
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 22369 4314 22435 4317
rect 26200 4314 27000 4344
rect 22369 4312 27000 4314
rect 22369 4256 22374 4312
rect 22430 4256 27000 4312
rect 22369 4254 27000 4256
rect 22369 4251 22435 4254
rect 26200 4224 27000 4254
rect 0 4178 800 4208
rect 3233 4178 3299 4181
rect 0 4176 3299 4178
rect 0 4120 3238 4176
rect 3294 4120 3299 4176
rect 0 4118 3299 4120
rect 0 4088 800 4118
rect 3233 4115 3299 4118
rect 7649 4178 7715 4181
rect 11646 4178 11652 4180
rect 7649 4176 11652 4178
rect 7649 4120 7654 4176
rect 7710 4120 11652 4176
rect 7649 4118 11652 4120
rect 7649 4115 7715 4118
rect 11646 4116 11652 4118
rect 11716 4116 11722 4180
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 8385 3770 8451 3773
rect 12566 3770 12572 3772
rect 8385 3768 12572 3770
rect 8385 3712 8390 3768
rect 8446 3712 12572 3768
rect 8385 3710 12572 3712
rect 8385 3707 8451 3710
rect 12566 3708 12572 3710
rect 12636 3708 12642 3772
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 5073 2954 5139 2957
rect 10542 2954 10548 2956
rect 5073 2952 10548 2954
rect 5073 2896 5078 2952
rect 5134 2896 10548 2952
rect 5073 2894 10548 2896
rect 5073 2891 5139 2894
rect 10542 2892 10548 2894
rect 10612 2892 10618 2956
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 14964 53892 15028 53956
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 14596 52592 14660 52596
rect 14596 52536 14610 52592
rect 14610 52536 14660 52592
rect 14596 52532 14660 52536
rect 22324 52532 22388 52596
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 17172 46412 17236 46476
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 15332 46004 15396 46068
rect 19748 45792 19812 45796
rect 19748 45736 19798 45792
rect 19798 45736 19812 45792
rect 19748 45732 19812 45736
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 19380 45596 19444 45660
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 20668 44780 20732 44844
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 10916 44236 10980 44300
rect 11836 44296 11900 44300
rect 11836 44240 11850 44296
rect 11850 44240 11900 44296
rect 11836 44236 11900 44240
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 12572 42876 12636 42940
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 21956 41516 22020 41580
rect 13676 41380 13740 41444
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 17724 40020 17788 40084
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 10916 38524 10980 38588
rect 12756 38524 12820 38588
rect 13676 38116 13740 38180
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 15148 37708 15212 37772
rect 17356 37708 17420 37772
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 20116 37300 20180 37364
rect 12572 37028 12636 37092
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 18644 36620 18708 36684
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 11836 36000 11900 36004
rect 11836 35944 11886 36000
rect 11886 35944 11900 36000
rect 11836 35940 11900 35944
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 12756 35124 12820 35188
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 12204 33764 12268 33828
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 17172 32540 17236 32604
rect 14596 32404 14660 32468
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 20116 31996 20180 32060
rect 15148 31724 15212 31788
rect 19932 31724 19996 31788
rect 22324 31724 22388 31788
rect 13676 31588 13740 31652
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 13492 30500 13556 30564
rect 24348 30560 24412 30564
rect 24348 30504 24398 30560
rect 24398 30504 24412 30560
rect 24348 30500 24412 30504
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 24532 30424 24596 30428
rect 24532 30368 24546 30424
rect 24546 30368 24596 30424
rect 24532 30364 24596 30368
rect 19380 30228 19444 30292
rect 19748 30228 19812 30292
rect 12572 30092 12636 30156
rect 15516 30092 15580 30156
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 17540 29472 17604 29476
rect 17540 29416 17590 29472
rect 17590 29416 17604 29472
rect 17540 29412 17604 29416
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 15516 29004 15580 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 14964 27508 15028 27572
rect 18460 27568 18524 27572
rect 18460 27512 18474 27568
rect 18474 27512 18524 27568
rect 18460 27508 18524 27512
rect 21956 27508 22020 27572
rect 20668 27372 20732 27436
rect 15332 27236 15396 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 14964 26828 15028 26892
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 14596 25060 14660 25124
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 15148 24924 15212 24988
rect 17172 24788 17236 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 17540 23488 17604 23492
rect 17540 23432 17590 23488
rect 17590 23432 17604 23488
rect 17540 23428 17604 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 11652 22476 11716 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 15516 21660 15580 21724
rect 13492 21524 13556 21588
rect 10548 21388 10612 21452
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 17356 20632 17420 20636
rect 17356 20576 17370 20632
rect 17370 20576 17420 20632
rect 17356 20572 17420 20576
rect 18644 20436 18708 20500
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18460 19348 18524 19412
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 20116 18804 20180 18868
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 12204 18396 12268 18460
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 15332 16552 15396 16556
rect 15332 16496 15382 16552
rect 15382 16496 15396 16552
rect 15332 16492 15396 16496
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 14964 16220 15028 16284
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 19932 15600 19996 15604
rect 19932 15544 19946 15600
rect 19946 15544 19996 15600
rect 19932 15540 19996 15544
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 24532 6760 24596 6764
rect 24532 6704 24546 6760
rect 24546 6704 24596 6760
rect 24532 6700 24596 6704
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 13492 5612 13556 5676
rect 24348 5612 24412 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 11652 4116 11716 4180
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 12572 3708 12636 3772
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 10548 2892 10612 2956
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 14963 53956 15029 53957
rect 14963 53892 14964 53956
rect 15028 53892 15029 53956
rect 14963 53891 15029 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 14595 52596 14661 52597
rect 14595 52532 14596 52596
rect 14660 52532 14661 52596
rect 14595 52531 14661 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 10915 44300 10981 44301
rect 10915 44236 10916 44300
rect 10980 44236 10981 44300
rect 10915 44235 10981 44236
rect 11835 44300 11901 44301
rect 11835 44236 11836 44300
rect 11900 44236 11901 44300
rect 11835 44235 11901 44236
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 10918 38589 10978 44235
rect 10915 38588 10981 38589
rect 10915 38524 10916 38588
rect 10980 38524 10981 38588
rect 10915 38523 10981 38524
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 11838 36005 11898 44235
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12571 42940 12637 42941
rect 12571 42876 12572 42940
rect 12636 42876 12637 42940
rect 12571 42875 12637 42876
rect 12574 37093 12634 42875
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 13675 41444 13741 41445
rect 13675 41380 13676 41444
rect 13740 41380 13741 41444
rect 13675 41379 13741 41380
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12755 38588 12821 38589
rect 12755 38524 12756 38588
rect 12820 38524 12821 38588
rect 12755 38523 12821 38524
rect 12571 37092 12637 37093
rect 12571 37028 12572 37092
rect 12636 37028 12637 37092
rect 12571 37027 12637 37028
rect 11835 36004 11901 36005
rect 11835 35940 11836 36004
rect 11900 35940 11901 36004
rect 11835 35939 11901 35940
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 12203 33828 12269 33829
rect 12203 33764 12204 33828
rect 12268 33764 12269 33828
rect 12203 33763 12269 33764
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 11651 22540 11717 22541
rect 11651 22476 11652 22540
rect 11716 22476 11717 22540
rect 11651 22475 11717 22476
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 10547 21452 10613 21453
rect 10547 21388 10548 21452
rect 10612 21388 10613 21452
rect 10547 21387 10613 21388
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 10550 2957 10610 21387
rect 11654 4181 11714 22475
rect 12206 18461 12266 33763
rect 12574 30157 12634 37027
rect 12758 35189 12818 38523
rect 12944 37568 13264 38592
rect 13678 38181 13738 41379
rect 13675 38180 13741 38181
rect 13675 38116 13676 38180
rect 13740 38116 13741 38180
rect 13675 38115 13741 38116
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12755 35188 12821 35189
rect 12755 35124 12756 35188
rect 12820 35124 12821 35188
rect 12755 35123 12821 35124
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 13678 31653 13738 38115
rect 14598 32469 14658 52531
rect 14595 32468 14661 32469
rect 14595 32404 14596 32468
rect 14660 32404 14661 32468
rect 14595 32403 14661 32404
rect 13675 31652 13741 31653
rect 13675 31588 13676 31652
rect 13740 31588 13741 31652
rect 13675 31587 13741 31588
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12571 30156 12637 30157
rect 12571 30092 12572 30156
rect 12636 30092 12637 30156
rect 12571 30091 12637 30092
rect 12203 18460 12269 18461
rect 12203 18396 12204 18460
rect 12268 18396 12269 18460
rect 12203 18395 12269 18396
rect 11651 4180 11717 4181
rect 11651 4116 11652 4180
rect 11716 4116 11717 4180
rect 11651 4115 11717 4116
rect 12574 3773 12634 30091
rect 12944 29952 13264 30976
rect 13491 30564 13557 30565
rect 13491 30500 13492 30564
rect 13556 30500 13557 30564
rect 13491 30499 13557 30500
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 13494 21589 13554 30499
rect 14598 25125 14658 32403
rect 14966 27573 15026 53891
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22323 52596 22389 52597
rect 22323 52532 22324 52596
rect 22388 52532 22389 52596
rect 22323 52531 22389 52532
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17171 46476 17237 46477
rect 17171 46412 17172 46476
rect 17236 46412 17237 46476
rect 17171 46411 17237 46412
rect 15331 46068 15397 46069
rect 15331 46004 15332 46068
rect 15396 46004 15397 46068
rect 15331 46003 15397 46004
rect 15147 37772 15213 37773
rect 15147 37708 15148 37772
rect 15212 37708 15213 37772
rect 15147 37707 15213 37708
rect 15150 31789 15210 37707
rect 15147 31788 15213 31789
rect 15147 31724 15148 31788
rect 15212 31724 15213 31788
rect 15147 31723 15213 31724
rect 15334 31770 15394 46003
rect 17174 32605 17234 46411
rect 17944 45728 18264 46752
rect 19747 45796 19813 45797
rect 19747 45732 19748 45796
rect 19812 45732 19813 45796
rect 19747 45731 19813 45732
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 19379 45660 19445 45661
rect 19379 45596 19380 45660
rect 19444 45596 19445 45660
rect 19379 45595 19445 45596
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17723 40084 17789 40085
rect 17723 40020 17724 40084
rect 17788 40020 17789 40084
rect 17723 40019 17789 40020
rect 17355 37772 17421 37773
rect 17355 37708 17356 37772
rect 17420 37708 17421 37772
rect 17355 37707 17421 37708
rect 17171 32604 17237 32605
rect 17171 32540 17172 32604
rect 17236 32540 17237 32604
rect 17171 32539 17237 32540
rect 14963 27572 15029 27573
rect 14963 27508 14964 27572
rect 15028 27508 15029 27572
rect 14963 27507 15029 27508
rect 14963 26892 15029 26893
rect 14963 26828 14964 26892
rect 15028 26828 15029 26892
rect 14963 26827 15029 26828
rect 14595 25124 14661 25125
rect 14595 25060 14596 25124
rect 14660 25060 14661 25124
rect 14595 25059 14661 25060
rect 13491 21588 13557 21589
rect 13491 21524 13492 21588
rect 13556 21524 13557 21588
rect 13491 21523 13557 21524
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 13494 5677 13554 21523
rect 14966 16285 15026 26827
rect 15150 24989 15210 31723
rect 15334 31710 15578 31770
rect 15518 30157 15578 31710
rect 15515 30156 15581 30157
rect 15515 30092 15516 30156
rect 15580 30092 15581 30156
rect 15515 30091 15581 30092
rect 15518 29069 15578 30091
rect 15515 29068 15581 29069
rect 15515 29004 15516 29068
rect 15580 29004 15581 29068
rect 15515 29003 15581 29004
rect 15331 27300 15397 27301
rect 15331 27236 15332 27300
rect 15396 27236 15397 27300
rect 15331 27235 15397 27236
rect 15147 24988 15213 24989
rect 15147 24924 15148 24988
rect 15212 24924 15213 24988
rect 15147 24923 15213 24924
rect 15334 16557 15394 27235
rect 15518 21725 15578 29003
rect 17174 24853 17234 32539
rect 17171 24852 17237 24853
rect 17171 24788 17172 24852
rect 17236 24788 17237 24852
rect 17171 24787 17237 24788
rect 15515 21724 15581 21725
rect 15515 21660 15516 21724
rect 15580 21660 15581 21724
rect 15515 21659 15581 21660
rect 17358 20637 17418 37707
rect 17726 31770 17786 40019
rect 17542 31710 17786 31770
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 18643 36684 18709 36685
rect 18643 36620 18644 36684
rect 18708 36620 18709 36684
rect 18643 36619 18709 36620
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17542 29477 17602 31710
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17539 29476 17605 29477
rect 17539 29412 17540 29476
rect 17604 29412 17605 29476
rect 17539 29411 17605 29412
rect 17542 23493 17602 29411
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 18459 27572 18525 27573
rect 18459 27508 18460 27572
rect 18524 27508 18525 27572
rect 18459 27507 18525 27508
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17539 23492 17605 23493
rect 17539 23428 17540 23492
rect 17604 23428 17605 23492
rect 17539 23427 17605 23428
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17355 20636 17421 20637
rect 17355 20572 17356 20636
rect 17420 20572 17421 20636
rect 17355 20571 17421 20572
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18462 19413 18522 27507
rect 18646 20501 18706 36619
rect 19382 30293 19442 45595
rect 19750 30293 19810 45731
rect 20667 44844 20733 44845
rect 20667 44780 20668 44844
rect 20732 44780 20733 44844
rect 20667 44779 20733 44780
rect 20115 37364 20181 37365
rect 20115 37300 20116 37364
rect 20180 37300 20181 37364
rect 20115 37299 20181 37300
rect 20118 32061 20178 37299
rect 20115 32060 20181 32061
rect 20115 31996 20116 32060
rect 20180 31996 20181 32060
rect 20115 31995 20181 31996
rect 19931 31788 19997 31789
rect 19931 31724 19932 31788
rect 19996 31724 19997 31788
rect 19931 31723 19997 31724
rect 19379 30292 19445 30293
rect 19379 30228 19380 30292
rect 19444 30228 19445 30292
rect 19379 30227 19445 30228
rect 19747 30292 19813 30293
rect 19747 30228 19748 30292
rect 19812 30228 19813 30292
rect 19747 30227 19813 30228
rect 18643 20500 18709 20501
rect 18643 20436 18644 20500
rect 18708 20436 18709 20500
rect 18643 20435 18709 20436
rect 18459 19412 18525 19413
rect 18459 19348 18460 19412
rect 18524 19348 18525 19412
rect 18459 19347 18525 19348
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 15331 16556 15397 16557
rect 15331 16492 15332 16556
rect 15396 16492 15397 16556
rect 15331 16491 15397 16492
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 14963 16284 15029 16285
rect 14963 16220 14964 16284
rect 15028 16220 15029 16284
rect 14963 16219 15029 16220
rect 17944 15264 18264 16288
rect 19934 15605 19994 31723
rect 20118 18869 20178 31995
rect 20670 27437 20730 44779
rect 21955 41580 22021 41581
rect 21955 41516 21956 41580
rect 22020 41516 22021 41580
rect 21955 41515 22021 41516
rect 21958 27573 22018 41515
rect 22326 31789 22386 52531
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22323 31788 22389 31789
rect 22323 31724 22324 31788
rect 22388 31724 22389 31788
rect 22323 31723 22389 31724
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 24347 30564 24413 30565
rect 24347 30500 24348 30564
rect 24412 30500 24413 30564
rect 24347 30499 24413 30500
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 21955 27572 22021 27573
rect 21955 27508 21956 27572
rect 22020 27508 22021 27572
rect 21955 27507 22021 27508
rect 20667 27436 20733 27437
rect 20667 27372 20668 27436
rect 20732 27372 20733 27436
rect 20667 27371 20733 27372
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 20115 18868 20181 18869
rect 20115 18804 20116 18868
rect 20180 18804 20181 18868
rect 20115 18803 20181 18804
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 19931 15604 19997 15605
rect 19931 15540 19932 15604
rect 19996 15540 19997 15604
rect 19931 15539 19997 15540
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 13491 5676 13557 5677
rect 13491 5612 13492 5676
rect 13556 5612 13557 5676
rect 13491 5611 13557 5612
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12571 3772 12637 3773
rect 12571 3708 12572 3772
rect 12636 3708 12637 3772
rect 12571 3707 12637 3708
rect 10547 2956 10613 2957
rect 10547 2892 10548 2956
rect 10612 2892 10613 2956
rect 10547 2891 10613 2892
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 24350 5677 24410 30499
rect 24531 30428 24597 30429
rect 24531 30364 24532 30428
rect 24596 30364 24597 30428
rect 24531 30363 24597 30364
rect 24534 6765 24594 30363
rect 24531 6764 24597 6765
rect 24531 6700 24532 6764
rect 24596 6700 24597 6764
rect 24531 6699 24597 6700
rect 24347 5676 24413 5677
rect 24347 5612 24348 5676
rect 24412 5612 24413 5676
rect 24347 5611 24413 5612
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_1  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1676037725
transform 1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _112_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 23828 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 23184 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 21160 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 23368 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 24104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 24840 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 24564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 16652 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 17848 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 18400 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 2668 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 3680 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 3864 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 6716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform 1 0 4140 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 4324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 5244 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1676037725
transform 1 0 6624 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 6256 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 6348 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 7084 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1676037725
transform 1 0 5888 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 7360 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 7544 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 8280 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform 1 0 6164 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 8464 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 8280 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 9660 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1676037725
transform 1 0 7820 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 10396 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 9936 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 11684 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 9292 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 9108 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform 1 0 12880 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 10488 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 11684 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 11776 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1676037725
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _206_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1676037725
transform 1 0 24564 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1676037725
transform 1 0 23736 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _209_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _210_
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _212_
timestamp 1676037725
transform 1 0 24564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 15548 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 17572 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 18676 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 20056 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3864 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4324 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8740 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6808 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8832 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10396 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6072 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5612 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5520 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13248 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13616 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12144 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10672 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7360 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__265 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12512 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__266
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4784 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 9936 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8096 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__267
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6992 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10304 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__268
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 8464 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6072 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3036 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3680 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 2852 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2576 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 2024 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 4416 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10212 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14536 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 20424 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 18124 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 11040 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 9016 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 11408 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 20516 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12
timestamp 1676037725
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1676037725
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1676037725
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1676037725
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1676037725
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1676037725
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_16
timestamp 1676037725
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1676037725
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1676037725
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1676037725
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_61
timestamp 1676037725
transform 1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1676037725
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_115
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1676037725
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1676037725
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1676037725
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_77
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_145
timestamp 1676037725
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1676037725
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1676037725
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_263
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_239
timestamp 1676037725
transform 1 0 23092 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_264
timestamp 1676037725
transform 1 0 25392 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1676037725
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1676037725
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_212
timestamp 1676037725
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_229
timestamp 1676037725
transform 1 0 22172 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1676037725
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1676037725
transform 1 0 19228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_202
timestamp 1676037725
transform 1 0 19688 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_212
timestamp 1676037725
transform 1 0 20608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_224
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1676037725
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_166
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_178
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1676037725
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1676037725
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1676037725
transform 1 0 14076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_146
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_242
timestamp 1676037725
transform 1 0 23368 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_117
timestamp 1676037725
transform 1 0 11868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1676037725
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1676037725
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1676037725
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1676037725
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_204
timestamp 1676037725
transform 1 0 19872 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_216
timestamp 1676037725
transform 1 0 20976 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1676037725
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1676037725
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1676037725
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1676037725
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_215
timestamp 1676037725
transform 1 0 20884 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_227
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_238
timestamp 1676037725
transform 1 0 23000 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_246
timestamp 1676037725
transform 1 0 23736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_195
timestamp 1676037725
transform 1 0 19044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1676037725
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_212
timestamp 1676037725
transform 1 0 20608 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_234
timestamp 1676037725
transform 1 0 22632 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1676037725
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_247
timestamp 1676037725
transform 1 0 23828 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1676037725
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_110
timestamp 1676037725
transform 1 0 11224 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1676037725
transform 1 0 12328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1676037725
transform 1 0 13064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_218
timestamp 1676037725
transform 1 0 21160 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_94
timestamp 1676037725
transform 1 0 9752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1676037725
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1676037725
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1676037725
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_117
timestamp 1676037725
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_127
timestamp 1676037725
transform 1 0 12788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_184
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_205
timestamp 1676037725
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1676037725
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1676037725
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1676037725
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1676037725
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1676037725
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 1676037725
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1676037725
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_207
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1676037725
transform 1 0 23644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1676037725
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_122
timestamp 1676037725
transform 1 0 12328 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_126
timestamp 1676037725
transform 1 0 12696 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1676037725
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1676037725
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_213
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_225
timestamp 1676037725
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_237
timestamp 1676037725
transform 1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1676037725
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_139
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1676037725
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_120
timestamp 1676037725
transform 1 0 12144 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1676037725
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_147
timestamp 1676037725
transform 1 0 14628 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_159
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_173
timestamp 1676037725
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1676037725
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 1676037725
transform 1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_100
timestamp 1676037725
transform 1 0 10304 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_197
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1676037725
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_254
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1676037725
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1676037725
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_72
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_78
timestamp 1676037725
transform 1 0 8280 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_96
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_162
timestamp 1676037725
transform 1 0 16008 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_174
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_229
timestamp 1676037725
transform 1 0 22172 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1676037725
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1676037725
transform 1 0 8280 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_91
timestamp 1676037725
transform 1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1676037725
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_141
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_151
timestamp 1676037725
transform 1 0 14996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1676037725
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1676037725
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_259
timestamp 1676037725
transform 1 0 24932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_37
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_60
timestamp 1676037725
transform 1 0 6624 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1676037725
transform 1 0 9660 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_108
timestamp 1676037725
transform 1 0 11040 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1676037725
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_219
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_231
timestamp 1676037725
transform 1 0 22356 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_83
timestamp 1676037725
transform 1 0 8740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1676037725
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_145
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 1676037725
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1676037725
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_202
timestamp 1676037725
transform 1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1676037725
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_255
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_263
timestamp 1676037725
transform 1 0 25300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_13
timestamp 1676037725
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1676037725
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_34
timestamp 1676037725
transform 1 0 4232 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_46
timestamp 1676037725
transform 1 0 5336 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1676037725
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1676037725
transform 1 0 10580 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_113
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1676037725
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1676037725
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_184
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1676037725
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1676037725
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1676037725
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1676037725
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_129
timestamp 1676037725
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1676037725
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1676037725
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_173
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_185
timestamp 1676037725
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1676037725
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1676037725
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1676037725
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_13
timestamp 1676037725
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1676037725
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_55
timestamp 1676037725
transform 1 0 6164 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_96
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_108
timestamp 1676037725
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 1676037725
transform 1 0 15916 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1676037725
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1676037725
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1676037725
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_232
timestamp 1676037725
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_77
timestamp 1676037725
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_102
timestamp 1676037725
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_124
timestamp 1676037725
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_136
timestamp 1676037725
transform 1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_180
timestamp 1676037725
transform 1 0 17664 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_212
timestamp 1676037725
transform 1 0 20608 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1676037725
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_51
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_63
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1676037725
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_126
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_202
timestamp 1676037725
transform 1 0 19688 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_23
timestamp 1676037725
transform 1 0 3220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_31
timestamp 1676037725
transform 1 0 3956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_35
timestamp 1676037725
transform 1 0 4324 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1676037725
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1676037725
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1676037725
transform 1 0 13524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1676037725
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1676037725
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_179
timestamp 1676037725
transform 1 0 17572 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_200
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1676037725
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_233
timestamp 1676037725
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_257
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1676037725
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1676037725
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1676037725
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1676037725
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_114
timestamp 1676037725
transform 1 0 11592 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_127
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_152
timestamp 1676037725
transform 1 0 15088 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_178
timestamp 1676037725
transform 1 0 17480 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_184
timestamp 1676037725
transform 1 0 18032 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1676037725
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_205
timestamp 1676037725
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_227
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_12
timestamp 1676037725
transform 1 0 2208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_24
timestamp 1676037725
transform 1 0 3312 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1676037725
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_80
timestamp 1676037725
transform 1 0 8464 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_104
timestamp 1676037725
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1676037725
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_153
timestamp 1676037725
transform 1 0 15180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1676037725
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_229
timestamp 1676037725
transform 1 0 22172 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1676037725
transform 1 0 22632 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_258
timestamp 1676037725
transform 1 0 24840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_47
timestamp 1676037725
transform 1 0 5428 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_68
timestamp 1676037725
transform 1 0 7360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1676037725
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_107
timestamp 1676037725
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_119
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1676037725
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_167
timestamp 1676037725
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1676037725
transform 1 0 17756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1676037725
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_217
timestamp 1676037725
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1676037725
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_77
timestamp 1676037725
transform 1 0 8188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_89
timestamp 1676037725
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1676037725
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1676037725
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_139
timestamp 1676037725
transform 1 0 13892 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_151
timestamp 1676037725
transform 1 0 14996 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1676037725
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1676037725
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1676037725
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_46
timestamp 1676037725
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_58
timestamp 1676037725
transform 1 0 6440 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_70
timestamp 1676037725
transform 1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_122
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1676037725
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1676037725
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_208
timestamp 1676037725
transform 1 0 20240 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_9
timestamp 1676037725
transform 1 0 1932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_13
timestamp 1676037725
transform 1 0 2300 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_41
timestamp 1676037725
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1676037725
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_70
timestamp 1676037725
transform 1 0 7544 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_94
timestamp 1676037725
transform 1 0 9752 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_100
timestamp 1676037725
transform 1 0 10304 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_136
timestamp 1676037725
transform 1 0 13616 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1676037725
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_192
timestamp 1676037725
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_265
timestamp 1676037725
transform 1 0 25484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_37
timestamp 1676037725
transform 1 0 4508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_49
timestamp 1676037725
transform 1 0 5612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_57
timestamp 1676037725
transform 1 0 6348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1676037725
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_90
timestamp 1676037725
transform 1 0 9384 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_98
timestamp 1676037725
transform 1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_105
timestamp 1676037725
transform 1 0 10764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_117
timestamp 1676037725
transform 1 0 11868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_129
timestamp 1676037725
transform 1 0 12972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1676037725
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_149
timestamp 1676037725
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_161
timestamp 1676037725
transform 1 0 15916 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_169
timestamp 1676037725
transform 1 0 16652 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1676037725
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_202
timestamp 1676037725
transform 1 0 19688 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_208
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_229
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_242
timestamp 1676037725
transform 1 0 23368 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_258
timestamp 1676037725
transform 1 0 24840 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_24
timestamp 1676037725
transform 1 0 3312 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_31
timestamp 1676037725
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_43
timestamp 1676037725
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_90
timestamp 1676037725
transform 1 0 9384 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_136
timestamp 1676037725
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_153
timestamp 1676037725
transform 1 0 15180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1676037725
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_186
timestamp 1676037725
transform 1 0 18216 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1676037725
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_211
timestamp 1676037725
transform 1 0 20516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_246
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_254
timestamp 1676037725
transform 1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_52
timestamp 1676037725
transform 1 0 5888 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_76
timestamp 1676037725
transform 1 0 8096 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_90
timestamp 1676037725
transform 1 0 9384 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_125
timestamp 1676037725
transform 1 0 12604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1676037725
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_212
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_220
timestamp 1676037725
transform 1 0 21344 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_242
timestamp 1676037725
transform 1 0 23368 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_13
timestamp 1676037725
transform 1 0 2300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_86
timestamp 1676037725
transform 1 0 9016 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_135
timestamp 1676037725
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_156
timestamp 1676037725
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_186
timestamp 1676037725
transform 1 0 18216 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp 1676037725
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_250
timestamp 1676037725
transform 1 0 24104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_254
timestamp 1676037725
transform 1 0 24472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_259
timestamp 1676037725
transform 1 0 24932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_265
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_52
timestamp 1676037725
transform 1 0 5888 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1676037725
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_106
timestamp 1676037725
transform 1 0 10856 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_118
timestamp 1676037725
transform 1 0 11960 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1676037725
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1676037725
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_156
timestamp 1676037725
transform 1 0 15456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1676037725
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1676037725
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_229
timestamp 1676037725
transform 1 0 22172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_259
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_79
timestamp 1676037725
transform 1 0 8372 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_87
timestamp 1676037725
transform 1 0 9108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1676037725
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_117
timestamp 1676037725
transform 1 0 11868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1676037725
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_142
timestamp 1676037725
transform 1 0 14168 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_152
timestamp 1676037725
transform 1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1676037725
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_208
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_240
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_244
timestamp 1676037725
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1676037725
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1676037725
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_52
timestamp 1676037725
transform 1 0 5888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_76
timestamp 1676037725
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_96
timestamp 1676037725
transform 1 0 9936 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_108
timestamp 1676037725
transform 1 0 11040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_130
timestamp 1676037725
transform 1 0 13064 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1676037725
transform 1 0 14444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_166
timestamp 1676037725
transform 1 0 16376 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_181
timestamp 1676037725
transform 1 0 17756 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_188
timestamp 1676037725
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_205
timestamp 1676037725
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_234
timestamp 1676037725
transform 1 0 22632 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_246
timestamp 1676037725
transform 1 0 23736 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_75
timestamp 1676037725
transform 1 0 8004 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_96
timestamp 1676037725
transform 1 0 9936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1676037725
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_145
timestamp 1676037725
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_213
timestamp 1676037725
transform 1 0 20700 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1676037725
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_230
timestamp 1676037725
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_242
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1676037725
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_259
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_265
timestamp 1676037725
transform 1 0 25484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_52
timestamp 1676037725
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_64
timestamp 1676037725
transform 1 0 6992 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_76
timestamp 1676037725
transform 1 0 8096 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_96
timestamp 1676037725
transform 1 0 9936 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_102
timestamp 1676037725
transform 1 0 10488 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_112
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_173
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1676037725
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1676037725
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_212
timestamp 1676037725
transform 1 0 20608 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_222
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_235
timestamp 1676037725
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1676037725
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_92
timestamp 1676037725
transform 1 0 9568 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_104
timestamp 1676037725
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_124
timestamp 1676037725
transform 1 0 12512 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_134
timestamp 1676037725
transform 1 0 13432 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_146
timestamp 1676037725
transform 1 0 14536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1676037725
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1676037725
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_180
timestamp 1676037725
transform 1 0 17664 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_188
timestamp 1676037725
transform 1 0 18400 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_206
timestamp 1676037725
transform 1 0 20056 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1676037725
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_61
timestamp 1676037725
transform 1 0 6716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_73
timestamp 1676037725
transform 1 0 7820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1676037725
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_163
timestamp 1676037725
transform 1 0 16100 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_171
timestamp 1676037725
transform 1 0 16836 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_182
timestamp 1676037725
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_229
timestamp 1676037725
transform 1 0 22172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1676037725
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_259
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_35
timestamp 1676037725
transform 1 0 4324 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_46
timestamp 1676037725
transform 1 0 5336 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1676037725
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_63
timestamp 1676037725
transform 1 0 6900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1676037725
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_80
timestamp 1676037725
transform 1 0 8464 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_92
timestamp 1676037725
transform 1 0 9568 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1676037725
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_175
timestamp 1676037725
transform 1 0 17204 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_185
timestamp 1676037725
transform 1 0 18124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_197
timestamp 1676037725
transform 1 0 19228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_209
timestamp 1676037725
transform 1 0 20332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_230
timestamp 1676037725
transform 1 0 22264 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_245
timestamp 1676037725
transform 1 0 23644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_253
timestamp 1676037725
transform 1 0 24380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_259
timestamp 1676037725
transform 1 0 24932 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_265
timestamp 1676037725
transform 1 0 25484 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_40
timestamp 1676037725
transform 1 0 4784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_64
timestamp 1676037725
transform 1 0 6992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_68
timestamp 1676037725
transform 1 0 7360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_78
timestamp 1676037725
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_107
timestamp 1676037725
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_119
timestamp 1676037725
transform 1 0 12052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1676037725
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_149
timestamp 1676037725
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_172
timestamp 1676037725
transform 1 0 16928 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_185
timestamp 1676037725
transform 1 0 18124 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1676037725
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_202
timestamp 1676037725
transform 1 0 19688 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_210
timestamp 1676037725
transform 1 0 20424 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_234
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_241
timestamp 1676037725
transform 1 0 23276 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_258
timestamp 1676037725
transform 1 0 24840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1676037725
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1676037725
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1676037725
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1676037725
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_72
timestamp 1676037725
transform 1 0 7728 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_83
timestamp 1676037725
transform 1 0 8740 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_108
timestamp 1676037725
transform 1 0 11040 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_131
timestamp 1676037725
transform 1 0 13156 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_135
timestamp 1676037725
transform 1 0 13524 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_143
timestamp 1676037725
transform 1 0 14260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1676037725
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_180
timestamp 1676037725
transform 1 0 17664 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_192
timestamp 1676037725
transform 1 0 18768 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_204
timestamp 1676037725
transform 1 0 19872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 1676037725
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1676037725
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1676037725
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_243
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_250
timestamp 1676037725
transform 1 0 24104 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_258
timestamp 1676037725
transform 1 0 24840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_47
timestamp 1676037725
transform 1 0 5428 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_68
timestamp 1676037725
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1676037725
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_96
timestamp 1676037725
transform 1 0 9936 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_108
timestamp 1676037725
transform 1 0 11040 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_114
timestamp 1676037725
transform 1 0 11592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_124
timestamp 1676037725
transform 1 0 12512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1676037725
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp 1676037725
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1676037725
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_191
timestamp 1676037725
transform 1 0 18676 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_203
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_229
timestamp 1676037725
transform 1 0 22172 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_242
timestamp 1676037725
transform 1 0 23368 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_246
timestamp 1676037725
transform 1 0 23736 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_92
timestamp 1676037725
transform 1 0 9568 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1676037725
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_143
timestamp 1676037725
transform 1 0 14260 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1676037725
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_194
timestamp 1676037725
transform 1 0 18952 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1676037725
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1676037725
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_61
timestamp 1676037725
transform 1 0 6716 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_73
timestamp 1676037725
transform 1 0 7820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1676037725
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_96
timestamp 1676037725
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_108
timestamp 1676037725
transform 1 0 11040 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_116
timestamp 1676037725
transform 1 0 11776 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1676037725
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_208
timestamp 1676037725
transform 1 0 20240 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_212
timestamp 1676037725
transform 1 0 20608 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1676037725
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1676037725
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_258
timestamp 1676037725
transform 1 0 24840 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1676037725
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_20
timestamp 1676037725
transform 1 0 2944 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1676037725
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1676037725
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_82
timestamp 1676037725
transform 1 0 8648 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_95
timestamp 1676037725
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1676037725
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_135
timestamp 1676037725
transform 1 0 13524 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_150
timestamp 1676037725
transform 1 0 14904 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_162
timestamp 1676037725
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_191
timestamp 1676037725
transform 1 0 18676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_204
timestamp 1676037725
transform 1 0 19872 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_211
timestamp 1676037725
transform 1 0 20516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1676037725
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_243
timestamp 1676037725
transform 1 0 23460 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_255
timestamp 1676037725
transform 1 0 24564 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1676037725
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_91
timestamp 1676037725
transform 1 0 9476 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_101
timestamp 1676037725
transform 1 0 10396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_113
timestamp 1676037725
transform 1 0 11500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_117
timestamp 1676037725
transform 1 0 11868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_158
timestamp 1676037725
transform 1 0 15640 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_170
timestamp 1676037725
transform 1 0 16744 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_182
timestamp 1676037725
transform 1 0 17848 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_214
timestamp 1676037725
transform 1 0 20792 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_226
timestamp 1676037725
transform 1 0 21896 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_234
timestamp 1676037725
transform 1 0 22632 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1676037725
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1676037725
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_136
timestamp 1676037725
transform 1 0 13616 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_162
timestamp 1676037725
transform 1 0 16008 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_180
timestamp 1676037725
transform 1 0 17664 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_188
timestamp 1676037725
transform 1 0 18400 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_210
timestamp 1676037725
transform 1 0 20424 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_74
timestamp 1676037725
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_98
timestamp 1676037725
transform 1 0 10120 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_106
timestamp 1676037725
transform 1 0 10856 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_119
timestamp 1676037725
transform 1 0 12052 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1676037725
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_156
timestamp 1676037725
transform 1 0 15456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_160
timestamp 1676037725
transform 1 0 15824 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_170
timestamp 1676037725
transform 1 0 16744 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_183
timestamp 1676037725
transform 1 0 17940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_214
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_220
timestamp 1676037725
transform 1 0 21344 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_230
timestamp 1676037725
transform 1 0 22264 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_238
timestamp 1676037725
transform 1 0 23000 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_8
timestamp 1676037725
transform 1 0 1840 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_20
timestamp 1676037725
transform 1 0 2944 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_32
timestamp 1676037725
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_90
timestamp 1676037725
transform 1 0 9384 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_103
timestamp 1676037725
transform 1 0 10580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_145
timestamp 1676037725
transform 1 0 14444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_150
timestamp 1676037725
transform 1 0 14904 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_163
timestamp 1676037725
transform 1 0 16100 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_174
timestamp 1676037725
transform 1 0 17112 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_182
timestamp 1676037725
transform 1 0 17848 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_201
timestamp 1676037725
transform 1 0 19596 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_211
timestamp 1676037725
transform 1 0 20516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1676037725
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_68
timestamp 1676037725
transform 1 0 7360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1676037725
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1676037725
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1676037725
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_120
timestamp 1676037725
transform 1 0 12144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_132
timestamp 1676037725
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_149
timestamp 1676037725
transform 1 0 14812 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_160
timestamp 1676037725
transform 1 0 15824 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1676037725
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1676037725
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_210
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_218
timestamp 1676037725
transform 1 0 21160 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_240
timestamp 1676037725
transform 1 0 23184 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1676037725
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1676037725
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1676037725
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_118
timestamp 1676037725
transform 1 0 11960 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_126
timestamp 1676037725
transform 1 0 12696 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_144
timestamp 1676037725
transform 1 0 14352 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_159
timestamp 1676037725
transform 1 0 15732 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_202
timestamp 1676037725
transform 1 0 19688 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_206
timestamp 1676037725
transform 1 0 20056 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_216
timestamp 1676037725
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_238
timestamp 1676037725
transform 1 0 23000 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_37
timestamp 1676037725
transform 1 0 4508 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_60
timestamp 1676037725
transform 1 0 6624 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_72
timestamp 1676037725
transform 1 0 7728 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1676037725
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_100
timestamp 1676037725
transform 1 0 10304 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_113
timestamp 1676037725
transform 1 0 11500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_117
timestamp 1676037725
transform 1 0 11868 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_127
timestamp 1676037725
transform 1 0 12788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_168
timestamp 1676037725
transform 1 0 16560 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_179
timestamp 1676037725
transform 1 0 17572 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_191
timestamp 1676037725
transform 1 0 18676 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_208
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_234
timestamp 1676037725
transform 1 0 22632 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_247
timestamp 1676037725
transform 1 0 23828 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_8
timestamp 1676037725
transform 1 0 1840 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_20
timestamp 1676037725
transform 1 0 2944 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_32
timestamp 1676037725
transform 1 0 4048 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_44
timestamp 1676037725
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_77
timestamp 1676037725
transform 1 0 8188 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_83
timestamp 1676037725
transform 1 0 8740 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_91
timestamp 1676037725
transform 1 0 9476 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_102
timestamp 1676037725
transform 1 0 10488 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1676037725
transform 1 0 11132 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_132
timestamp 1676037725
transform 1 0 13248 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_145
timestamp 1676037725
transform 1 0 14444 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_153
timestamp 1676037725
transform 1 0 15180 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1676037725
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_177
timestamp 1676037725
transform 1 0 17388 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_200
timestamp 1676037725
transform 1 0 19504 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_213
timestamp 1676037725
transform 1 0 20700 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1676037725
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_236
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_263
timestamp 1676037725
transform 1 0 25300 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_80
timestamp 1676037725
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_96
timestamp 1676037725
transform 1 0 9936 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_134
timestamp 1676037725
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_152
timestamp 1676037725
transform 1 0 15088 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_158
timestamp 1676037725
transform 1 0 15640 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_168
timestamp 1676037725
transform 1 0 16560 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_176
timestamp 1676037725
transform 1 0 17296 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_186
timestamp 1676037725
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_222
timestamp 1676037725
transform 1 0 21528 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_235
timestamp 1676037725
transform 1 0 22724 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1676037725
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_82
timestamp 1676037725
transform 1 0 8648 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_97
timestamp 1676037725
transform 1 0 10028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_109
timestamp 1676037725
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_119
timestamp 1676037725
transform 1 0 12052 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_140
timestamp 1676037725
transform 1 0 13984 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_147
timestamp 1676037725
transform 1 0 14628 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_162
timestamp 1676037725
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_236
timestamp 1676037725
transform 1 0 22816 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_250
timestamp 1676037725
transform 1 0 24104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_76
timestamp 1676037725
transform 1 0 8096 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_123
timestamp 1676037725
transform 1 0 12420 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_136
timestamp 1676037725
transform 1 0 13616 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_159
timestamp 1676037725
transform 1 0 15732 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_169
timestamp 1676037725
transform 1 0 16652 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_175
timestamp 1676037725
transform 1 0 17204 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_185
timestamp 1676037725
transform 1 0 18124 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_193
timestamp 1676037725
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_208
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_216
timestamp 1676037725
transform 1 0 20976 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_237
timestamp 1676037725
transform 1 0 22908 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_258
timestamp 1676037725
transform 1 0 24840 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_34
timestamp 1676037725
transform 1 0 4232 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_46
timestamp 1676037725
transform 1 0 5336 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1676037725
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_79
timestamp 1676037725
transform 1 0 8372 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_87
timestamp 1676037725
transform 1 0 9108 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1676037725
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_124
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_132
timestamp 1676037725
transform 1 0 13248 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_153
timestamp 1676037725
transform 1 0 15180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_165
timestamp 1676037725
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_180
timestamp 1676037725
transform 1 0 17664 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_71_208
timestamp 1676037725
transform 1 0 20240 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_216
timestamp 1676037725
transform 1 0 20976 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1676037725
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_260
timestamp 1676037725
transform 1 0 25024 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_9
timestamp 1676037725
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_39
timestamp 1676037725
transform 1 0 4692 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_49
timestamp 1676037725
transform 1 0 5612 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_61
timestamp 1676037725
transform 1 0 6716 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_82
timestamp 1676037725
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_174
timestamp 1676037725
transform 1 0 17112 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_182
timestamp 1676037725
transform 1 0 17848 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_208
timestamp 1676037725
transform 1 0 20240 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_220
timestamp 1676037725
transform 1 0 21344 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_231
timestamp 1676037725
transform 1 0 22356 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_239
timestamp 1676037725
transform 1 0 23092 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_32
timestamp 1676037725
transform 1 0 4048 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_44
timestamp 1676037725
transform 1 0 5152 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_124
timestamp 1676037725
transform 1 0 12512 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_156
timestamp 1676037725
transform 1 0 15456 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_202
timestamp 1676037725
transform 1 0 19688 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_210
timestamp 1676037725
transform 1 0 20424 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_236
timestamp 1676037725
transform 1 0 22816 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_240
timestamp 1676037725
transform 1 0 23184 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_265
timestamp 1676037725
transform 1 0 25484 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_37
timestamp 1676037725
transform 1 0 4508 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_49
timestamp 1676037725
transform 1 0 5612 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_55
timestamp 1676037725
transform 1 0 6164 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_60
timestamp 1676037725
transform 1 0 6624 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_67
timestamp 1676037725
transform 1 0 7268 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_74
timestamp 1676037725
transform 1 0 7912 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1676037725
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_89
timestamp 1676037725
transform 1 0 9292 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_99
timestamp 1676037725
transform 1 0 10212 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_111
timestamp 1676037725
transform 1 0 11316 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_117
timestamp 1676037725
transform 1 0 11868 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_127
timestamp 1676037725
transform 1 0 12788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_163
timestamp 1676037725
transform 1 0 16100 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_175
timestamp 1676037725
transform 1 0 17204 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_187
timestamp 1676037725
transform 1 0 18308 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_219
timestamp 1676037725
transform 1 0 21252 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_227
timestamp 1676037725
transform 1 0 21988 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1676037725
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_47
timestamp 1676037725
transform 1 0 5428 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_102
timestamp 1676037725
transform 1 0 10488 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1676037725
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_130
timestamp 1676037725
transform 1 0 13064 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_142
timestamp 1676037725
transform 1 0 14168 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_154
timestamp 1676037725
transform 1 0 15272 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_180
timestamp 1676037725
transform 1 0 17664 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_192
timestamp 1676037725
transform 1 0 18768 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_204
timestamp 1676037725
transform 1 0 19872 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_216
timestamp 1676037725
transform 1 0 20976 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_247
timestamp 1676037725
transform 1 0 23828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_253
timestamp 1676037725
transform 1 0 24380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_61
timestamp 1676037725
transform 1 0 6716 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_73
timestamp 1676037725
transform 1 0 7820 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1676037725
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_105
timestamp 1676037725
transform 1 0 10764 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_113
timestamp 1676037725
transform 1 0 11500 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1676037725
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_159
timestamp 1676037725
transform 1 0 15732 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_180
timestamp 1676037725
transform 1 0 17664 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_192
timestamp 1676037725
transform 1 0 18768 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_219
timestamp 1676037725
transform 1 0 21252 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_227
timestamp 1676037725
transform 1 0 21988 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_249
timestamp 1676037725
transform 1 0 24012 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_264
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_76
timestamp 1676037725
transform 1 0 8096 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_84
timestamp 1676037725
transform 1 0 8832 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1676037725
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_124
timestamp 1676037725
transform 1 0 12512 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_132
timestamp 1676037725
transform 1 0 13248 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_140
timestamp 1676037725
transform 1 0 13984 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1676037725
transform 1 0 16100 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_177
timestamp 1676037725
transform 1 0 17388 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_200
timestamp 1676037725
transform 1 0 19504 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_212
timestamp 1676037725
transform 1 0 20608 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_77_247
timestamp 1676037725
transform 1 0 23828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_253
timestamp 1676037725
transform 1 0 24380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_257
timestamp 1676037725
transform 1 0 24748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_72
timestamp 1676037725
transform 1 0 7728 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_93
timestamp 1676037725
transform 1 0 9660 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_100
timestamp 1676037725
transform 1 0 10304 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_124
timestamp 1676037725
transform 1 0 12512 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_136
timestamp 1676037725
transform 1 0 13616 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_163
timestamp 1676037725
transform 1 0 16100 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_175
timestamp 1676037725
transform 1 0 17204 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_187
timestamp 1676037725
transform 1 0 18308 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_219
timestamp 1676037725
transform 1 0 21252 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_232
timestamp 1676037725
transform 1 0 22448 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_258
timestamp 1676037725
transform 1 0 24840 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_77
timestamp 1676037725
transform 1 0 8188 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_82
timestamp 1676037725
transform 1 0 8648 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_97
timestamp 1676037725
transform 1 0 10028 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_110
timestamp 1676037725
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_119
timestamp 1676037725
transform 1 0 12052 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_131
timestamp 1676037725
transform 1 0 13156 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_153
timestamp 1676037725
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1676037725
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_191
timestamp 1676037725
transform 1 0 18676 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_199
timestamp 1676037725
transform 1 0 19412 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_211
timestamp 1676037725
transform 1 0 20516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_245
timestamp 1676037725
transform 1 0 23644 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_69
timestamp 1676037725
transform 1 0 7452 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_74
timestamp 1676037725
transform 1 0 7912 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_159
timestamp 1676037725
transform 1 0 15732 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_180
timestamp 1676037725
transform 1 0 17664 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_192
timestamp 1676037725
transform 1 0 18768 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_208
timestamp 1676037725
transform 1 0 20240 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_223
timestamp 1676037725
transform 1 0 21620 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_235
timestamp 1676037725
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1676037725
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_63
timestamp 1676037725
transform 1 0 6900 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_67
timestamp 1676037725
transform 1 0 7268 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_79
timestamp 1676037725
transform 1 0 8372 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_91
timestamp 1676037725
transform 1 0 9476 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_103
timestamp 1676037725
transform 1 0 10580 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_133
timestamp 1676037725
transform 1 0 13340 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_156
timestamp 1676037725
transform 1 0 15456 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_180
timestamp 1676037725
transform 1 0 17664 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_265
timestamp 1676037725
transform 1 0 25484 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_90
timestamp 1676037725
transform 1 0 9384 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_102
timestamp 1676037725
transform 1 0 10488 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_110
timestamp 1676037725
transform 1 0 11224 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_116
timestamp 1676037725
transform 1 0 11776 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_128
timestamp 1676037725
transform 1 0 12880 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_149
timestamp 1676037725
transform 1 0 14812 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_172
timestamp 1676037725
transform 1 0 16928 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_185
timestamp 1676037725
transform 1 0 18124 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1676037725
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_257
timestamp 1676037725
transform 1 0 24748 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_54
timestamp 1676037725
transform 1 0 6072 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_118
timestamp 1676037725
transform 1 0 11960 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_130
timestamp 1676037725
transform 1 0 13064 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_142
timestamp 1676037725
transform 1 0 14168 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_154
timestamp 1676037725
transform 1 0 15272 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_166
timestamp 1676037725
transform 1 0 16376 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_257
timestamp 1676037725
transform 1 0 24748 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_264
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_259
timestamp 1676037725
transform 1 0 24932 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_23
timestamp 1676037725
transform 1 0 3220 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_35
timestamp 1676037725
transform 1 0 4324 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_47
timestamp 1676037725
transform 1 0 5428 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_76
timestamp 1676037725
transform 1 0 8096 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_88
timestamp 1676037725
transform 1 0 9200 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_265
timestamp 1676037725
transform 1 0 25484 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1676037725
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_47
timestamp 1676037725
transform 1 0 5428 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_58
timestamp 1676037725
transform 1 0 6440 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_70
timestamp 1676037725
transform 1 0 7544 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_82
timestamp 1676037725
transform 1 0 8648 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1676037725
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1676037725
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1676037725
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1676037725
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_259
timestamp 1676037725
transform 1 0 24932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_264
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_35
timestamp 1676037725
transform 1 0 4324 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_47
timestamp 1676037725
transform 1 0 5428 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_65
timestamp 1676037725
transform 1 0 7084 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_77
timestamp 1676037725
transform 1 0 8188 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_89
timestamp 1676037725
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_97
timestamp 1676037725
transform 1 0 10028 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_101
timestamp 1676037725
transform 1 0 10396 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_257
timestamp 1676037725
transform 1 0 24748 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1676037725
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_47
timestamp 1676037725
transform 1 0 5428 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_51
timestamp 1676037725
transform 1 0 5796 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_55
timestamp 1676037725
transform 1 0 6164 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_75
timestamp 1676037725
transform 1 0 8004 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_259
timestamp 1676037725
transform 1 0 24932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1676037725
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1676037725
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_79
timestamp 1676037725
transform 1 0 8372 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1676037725
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_118
timestamp 1676037725
transform 1 0 11960 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_130
timestamp 1676037725
transform 1 0 13064 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_142
timestamp 1676037725
transform 1 0 14168 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_154
timestamp 1676037725
transform 1 0 15272 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_166
timestamp 1676037725
transform 1 0 16376 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_257
timestamp 1676037725
transform 1 0 24748 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1676037725
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1676037725
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1676037725
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_93
timestamp 1676037725
transform 1 0 9660 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_111
timestamp 1676037725
transform 1 0 11316 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_115
timestamp 1676037725
transform 1 0 11684 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_119
timestamp 1676037725
transform 1 0 12052 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_126
timestamp 1676037725
transform 1 0 12696 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_130
timestamp 1676037725
transform 1 0 13064 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_135
timestamp 1676037725
transform 1 0 13524 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_249
timestamp 1676037725
transform 1 0 24012 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_8
timestamp 1676037725
transform 1 0 1840 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_16
timestamp 1676037725
transform 1 0 2576 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1676037725
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_93_63
timestamp 1676037725
transform 1 0 6900 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_71
timestamp 1676037725
transform 1 0 7636 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1676037725
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_131
timestamp 1676037725
transform 1 0 13156 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_139
timestamp 1676037725
transform 1 0 13892 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_147
timestamp 1676037725
transform 1 0 14628 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_159
timestamp 1676037725
transform 1 0 15732 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_201
timestamp 1676037725
transform 1 0 19596 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_206
timestamp 1676037725
transform 1 0 20056 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_218
timestamp 1676037725
transform 1 0 21160 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_231
timestamp 1676037725
transform 1 0 22356 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_238
timestamp 1676037725
transform 1 0 23000 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_246
timestamp 1676037725
transform 1 0 23736 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1676037725
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_111
timestamp 1676037725
transform 1 0 11316 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_131
timestamp 1676037725
transform 1 0 13156 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_138
timestamp 1676037725
transform 1 0 13800 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_147
timestamp 1676037725
transform 1 0 14628 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_163
timestamp 1676037725
transform 1 0 16100 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_171
timestamp 1676037725
transform 1 0 16836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_178
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_182
timestamp 1676037725
transform 1 0 17848 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_187
timestamp 1676037725
transform 1 0 18308 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_203
timestamp 1676037725
transform 1 0 19780 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_223
timestamp 1676037725
transform 1 0 21620 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_230
timestamp 1676037725
transform 1 0 22264 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_258
timestamp 1676037725
transform 1 0 24840 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_135
timestamp 1676037725
transform 1 0 13524 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_139
timestamp 1676037725
transform 1 0 13892 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_151
timestamp 1676037725
transform 1 0 14996 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_159
timestamp 1676037725
transform 1 0 15732 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1676037725
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_191
timestamp 1676037725
transform 1 0 18676 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1676037725
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1676037725
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1676037725
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_219
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_230
timestamp 1676037725
transform 1 0 22264 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_258
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 23552 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 25116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 24472 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 23184 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 23184 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 24472 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 24472 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23276 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1676037725
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1676037725
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 12420 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 16468 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17204 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 17940 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 18676 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 19412 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 20148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 14260 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 19780 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 20884 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 20516 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21252 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 21988 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 22724 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 13156 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform 1 0 13524 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 13524 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform 1 0 14260 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 14628 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 15364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 16100 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 15732 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1676037725
transform 1 0 25024 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1676037725
transform 1 0 25024 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 25024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 25024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1676037725
transform 1 0 25024 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input108
timestamp 1676037725
transform 1 0 22264 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112
timestamp 1676037725
transform 1 0 3956 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  left_tile_264
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output113 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 3956 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 22080 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 22080 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 23920 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 22080 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 23920 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 4600 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 5336 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 6532 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 6900 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 7176 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 1748 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 7912 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 9108 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 9844 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 9844 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 11684 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 11684 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2024 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 2024 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 2852 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 2024 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 2760 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 3956 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 2760 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output211
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output212
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output213
timestamp 1676037725
transform 1 0 23920 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output214
timestamp 1676037725
transform 1 0 22632 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output215
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output216
timestamp 1676037725
transform 1 0 23920 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output217
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output218
timestamp 1676037725
transform 1 0 22632 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23000 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22632 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20148 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19596 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14536 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19320 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23276 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22172 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14536 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15088 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14444 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20700 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23184 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21068 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21344 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22724 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23184 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23552 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22172 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18400 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17848 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17664 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15824 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15824 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15088 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13616 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13616 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11960 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10764 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11224 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8096 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6256 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6256 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6256 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6440 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7912 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8832 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11224 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14996 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22724 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 -1 48960
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10672 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12144 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9384 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10304 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7544 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7544 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6072 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4784 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5244 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5244 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6716 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7728 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 7728 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5152 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 5520 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 3496 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4232 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6256 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7820 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11316 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15272 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17664 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17020 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__269
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14352 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21896 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20608 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 20792 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22908 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20424 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16928 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__224
timestamp 1676037725
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19044 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15548 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__270
timestamp 1676037725
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15456 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20516 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__271
timestamp 1676037725
transform 1 0 20240 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19136 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22540 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19780 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__272
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19964 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__273
timestamp 1676037725
transform 1 0 18124 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16928 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 13156 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12696 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__223
timestamp 1676037725
transform 1 0 14628 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15272 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11316 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21804 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__225
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21804 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23920 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21804 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20608 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21896 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__242
timestamp 1676037725
transform 1 0 20240 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19044 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23368 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21528 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23000 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__251
timestamp 1676037725
transform 1 0 23184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22816 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20700 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 21252 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19504 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__226
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15916 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__227
timestamp 1676037725
transform 1 0 19412 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16376 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15732 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__228
timestamp 1676037725
transform 1 0 16100 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 14352 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13616 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19504 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__230
timestamp 1676037725
transform 1 0 14076 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12880 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14168 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12880 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 13248 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14628 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19136 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12788 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13432 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14628 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__234
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12144 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__235
timestamp 1676037725
transform 1 0 10580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10120 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 8740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7544 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__237
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 7268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__239
timestamp 1676037725
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__240
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8924 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__243
timestamp 1676037725
transform 1 0 16652 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__244
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__246
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__247
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 23092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9384 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17296 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15180 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__253
timestamp 1676037725
transform 1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 10120 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11868 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__256
timestamp 1676037725
transform 1 0 12972 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11776 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14352 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18124 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 10120 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12880 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 10948 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9568 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12972 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__263
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 6992 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9476 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9016 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7820 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__254
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 6992 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9752 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9936 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7728 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7820 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13984 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17296 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__255
timestamp 1676037725
transform 1 0 8464 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9752 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7636 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14076 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7452 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__257
timestamp 1676037725
transform 1 0 8188 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6992 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12420 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12328 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__258
timestamp 1676037725
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 4508 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5152 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5520 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__259
timestamp 1676037725
transform 1 0 8464 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6992 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10672 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__261
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19688 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14812 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 4224 27000 4344 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 938 56200 994 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25304 27000 25424 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 32104 27000 32224 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 32784 27000 32904 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 33464 27000 33584 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 34824 27000 34944 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 35504 27000 35624 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 36184 27000 36304 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 36864 27000 36984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 37544 27000 37664 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 38904 27000 39024 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 39584 27000 39704 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 40264 27000 40384 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 40944 27000 41064 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 41624 27000 41744 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 42984 27000 43104 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 43664 27000 43784 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 44344 27000 44464 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 45024 27000 45144 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 26664 27000 26784 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 27344 27000 27464 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 28024 27000 28144 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 28704 27000 28824 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 29384 27000 29504 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 30744 27000 30864 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 31424 27000 31544 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 4904 27000 5024 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 12384 27000 12504 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 13064 27000 13184 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 14424 27000 14544 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 15104 27000 15224 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 16464 27000 16584 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 17144 27000 17264 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 18504 27000 18624 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 19184 27000 19304 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20544 27000 20664 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21224 27000 21344 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22584 27000 22704 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23264 27000 23384 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 24624 27000 24744 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 6264 27000 6384 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 6944 27000 7064 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 8304 27000 8424 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 8984 27000 9104 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 10344 27000 10464 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 11024 27000 11144 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12346 56200 12402 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16026 56200 16082 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16394 56200 16450 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 16762 56200 16818 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17130 56200 17186 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 17498 56200 17554 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 17866 56200 17922 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18234 56200 18290 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 18602 56200 18658 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19338 56200 19394 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 12714 56200 12770 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 19706 56200 19762 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20074 56200 20130 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20442 56200 20498 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 20810 56200 20866 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21178 56200 21234 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 21546 56200 21602 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 21914 56200 21970 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22282 56200 22338 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 22650 56200 22706 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23018 56200 23074 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13082 56200 13138 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 13818 56200 13874 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14186 56200 14242 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 14554 56200 14610 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 14922 56200 14978 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15290 56200 15346 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 15658 56200 15714 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1306 56200 1362 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 4986 56200 5042 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5354 56200 5410 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 5722 56200 5778 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6090 56200 6146 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 6458 56200 6514 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 6826 56200 6882 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7194 56200 7250 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 7562 56200 7618 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8298 56200 8354 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 1674 56200 1730 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 8666 56200 8722 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9034 56200 9090 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9402 56200 9458 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 9770 56200 9826 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10138 56200 10194 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 10506 56200 10562 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 10874 56200 10930 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11242 56200 11298 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 11610 56200 11666 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 11978 56200 12034 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2042 56200 2098 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 2778 56200 2834 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3146 56200 3202 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 3514 56200 3570 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 3882 56200 3938 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4250 56200 4306 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 4618 56200 4674 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 36456 800 36576 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 24896 800 25016 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 200 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_reset_bottom_out
port 201 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 prog_reset_left_in
port 202 nsew signal input
flabel metal3 s 26200 45704 27000 45824 0 FreeSans 480 0 0 0 prog_reset_right_out
port 203 nsew signal tristate
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 204 nsew signal input
flabel metal2 s 24122 56200 24178 57000 0 FreeSans 224 90 0 0 prog_reset_top_out
port 205 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 206 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset_bottom_out
port 207 nsew signal tristate
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 reset_right_in
port 208 nsew signal input
flabel metal2 s 25226 56200 25282 57000 0 FreeSans 224 90 0 0 reset_top_in
port 209 nsew signal input
flabel metal2 s 24858 56200 24914 57000 0 FreeSans 224 90 0 0 reset_top_out
port 210 nsew signal tristate
flabel metal3 s 26200 47064 27000 47184 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 211 nsew signal input
flabel metal3 s 26200 47744 27000 47864 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 212 nsew signal input
flabel metal3 s 26200 48424 27000 48544 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 213 nsew signal input
flabel metal3 s 26200 49104 27000 49224 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 214 nsew signal input
flabel metal3 s 26200 49784 27000 49904 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 215 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 216 nsew signal input
flabel metal3 s 26200 51144 27000 51264 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 217 nsew signal input
flabel metal3 s 26200 51824 27000 51944 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 218 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 219 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 220 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 221 nsew signal tristate
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 222 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 223 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 test_enable_bottom_out
port 224 nsew signal tristate
flabel metal3 s 26200 52504 27000 52624 0 FreeSans 480 0 0 0 test_enable_right_in
port 225 nsew signal input
flabel metal2 s 25962 56200 26018 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 226 nsew signal input
flabel metal2 s 25594 56200 25650 57000 0 FreeSans 224 90 0 0 test_enable_top_out
port 227 nsew signal tristate
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 228 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 229 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 230 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 231 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal2 6026 24276 6026 24276 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 3726 23290 3726 23290 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 3726 22474 3726 22474 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 3910 18938 3910 18938 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 2806 21148 2806 21148 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7038 19890 7038 19890 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 9338 8534 9338 8534 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal2 7958 20077 7958 20077 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 7820 22134 7820 22134 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 8602 14110 8602 14110 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 11960 22134 11960 22134 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13248 14926 13248 14926 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 10442 14790 10442 14790 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6256 17102 6256 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 15502 11186 15502 11186 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 12282 14246 12282 14246 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 7452 16014 7452 16014 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal2 12236 22508 12236 22508 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 10350 20774 10350 20774 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal2 5842 23392 5842 23392 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 12742 15538 12742 15538 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7314 21760 7314 21760 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 5014 23018 5014 23018 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13294 17068 13294 17068 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12190 19244 12190 19244 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12144 20570 12144 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9660 18938 9660 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 10166 18496 10166 18496 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10074 19822 10074 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7590 20570 7590 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8602 21998 8602 21998 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 9154 20808 9154 20808 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 14950 12138 14950 12138 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8556 15130 8556 15130 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 7590 17238 7590 17238 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14168 15130 14168 15130 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 17646 13662 17646 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13616 17578 13616 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10764 21862 10764 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12972 15130 12972 15130 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12558 16966 12558 16966 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9430 14586 9430 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10212 16558 10212 16558 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7958 15062 7958 15062 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15502 11016 15502 11016 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7038 16694 7038 16694 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4738 17306 4738 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13938 11254 13938 11254 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12604 17238 12604 17238 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12098 17952 12098 17952 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9154 19482 9154 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11776 12954 11776 12954 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10856 16966 10856 16966 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7498 17850 7498 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8786 16014 8786 16014 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 7222 17306 7222 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 11822 17000 11822 17000 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 5888 22202 5888 22202 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4738 22406 4738 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 11730 18870 11730 18870 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11638 20128 11638 20128 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11132 20910 11132 20910 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8970 16422 8970 16422 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10350 19482 10350 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9246 21114 9246 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7130 21114 7130 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7498 21930 7498 21930 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6716 22610 6716 22610 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4738 24582 4738 24582 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 3220 25806 3220 25806 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 2944 25738 2944 25738 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel via1 3519 27098 3519 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4048 23494 4048 23494 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 3404 24038 3404 24038 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 3082 22746 3082 22746 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 3933 26010 3933 26010 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 5750 18224 5750 18224 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 2484 21454 2484 21454 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 2944 22100 2944 22100 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel via1 4117 24378 4117 24378 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 3743 22610 3743 22610 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 3036 21114 3036 21114 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 3979 22746 3979 22746 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 1740 55012 1740 55012 0 ccff_head
rlabel metal3 1740 1836 1740 1836 0 ccff_head_0
rlabel metal1 21850 6358 21850 6358 0 ccff_tail
rlabel metal1 2714 52598 2714 52598 0 ccff_tail_0
rlabel metal2 22310 25619 22310 25619 0 chanx_right_in[0]
rlabel metal2 25346 32521 25346 32521 0 chanx_right_in[10]
rlabel metal1 24472 32878 24472 32878 0 chanx_right_in[11]
rlabel metal2 25346 34051 25346 34051 0 chanx_right_in[12]
rlabel metal1 25392 35054 25392 35054 0 chanx_right_in[13]
rlabel metal1 25438 36142 25438 36142 0 chanx_right_in[14]
rlabel metal2 25346 36159 25346 36159 0 chanx_right_in[15]
rlabel metal1 25392 38318 25392 38318 0 chanx_right_in[16]
rlabel metal1 24840 37230 24840 37230 0 chanx_right_in[17]
rlabel metal2 23782 37417 23782 37417 0 chanx_right_in[18]
rlabel metal3 25860 38284 25860 38284 0 chanx_right_in[19]
rlabel metal1 25070 24174 25070 24174 0 chanx_right_in[1]
rlabel metal1 24518 39916 24518 39916 0 chanx_right_in[20]
rlabel metal1 24058 40018 24058 40018 0 chanx_right_in[21]
rlabel metal2 24058 39865 24058 39865 0 chanx_right_in[22]
rlabel metal3 24802 41004 24802 41004 0 chanx_right_in[23]
rlabel metal2 25346 42177 25346 42177 0 chanx_right_in[24]
rlabel metal1 25070 43758 25070 43758 0 chanx_right_in[25]
rlabel metal1 24702 43282 24702 43282 0 chanx_right_in[26]
rlabel metal2 25346 44047 25346 44047 0 chanx_right_in[27]
rlabel metal1 24794 44370 24794 44370 0 chanx_right_in[28]
rlabel metal3 25538 45084 25538 45084 0 chanx_right_in[29]
rlabel metal2 23506 27387 23506 27387 0 chanx_right_in[2]
rlabel metal1 24518 26350 24518 26350 0 chanx_right_in[3]
rlabel metal1 24472 28526 24472 28526 0 chanx_right_in[4]
rlabel metal2 24150 28951 24150 28951 0 chanx_right_in[5]
rlabel metal2 25346 28985 25346 28985 0 chanx_right_in[6]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[7]
rlabel metal1 25392 32402 25392 32402 0 chanx_right_in[8]
rlabel metal3 25216 31484 25216 31484 0 chanx_right_in[9]
rlabel metal3 25860 11764 25860 11764 0 chanx_right_out[10]
rlabel metal1 24104 12886 24104 12886 0 chanx_right_out[11]
rlabel metal2 24702 12393 24702 12393 0 chanx_right_out[12]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[13]
rlabel metal1 24104 15062 24104 15062 0 chanx_right_out[14]
rlabel metal2 25162 14569 25162 14569 0 chanx_right_out[15]
rlabel metal1 24380 15538 24380 15538 0 chanx_right_out[16]
rlabel metal2 24794 15725 24794 15725 0 chanx_right_out[17]
rlabel metal3 25124 17204 25124 17204 0 chanx_right_out[18]
rlabel metal1 22310 18088 22310 18088 0 chanx_right_out[19]
rlabel metal2 24794 5389 24794 5389 0 chanx_right_out[1]
rlabel metal2 23874 18139 23874 18139 0 chanx_right_out[20]
rlabel metal2 22218 19329 22218 19329 0 chanx_right_out[21]
rlabel metal1 24104 19414 24104 19414 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel metal2 24702 20281 24702 20281 0 chanx_right_out[24]
rlabel metal3 25676 21964 25676 21964 0 chanx_right_out[25]
rlabel metal3 26228 22644 26228 22644 0 chanx_right_out[26]
rlabel metal1 23368 23630 23368 23630 0 chanx_right_out[27]
rlabel metal3 25676 24004 25676 24004 0 chanx_right_out[28]
rlabel metal2 25162 24225 25162 24225 0 chanx_right_out[29]
rlabel metal3 25676 6324 25676 6324 0 chanx_right_out[2]
rlabel metal3 25584 7004 25584 7004 0 chanx_right_out[3]
rlabel metal3 25676 7684 25676 7684 0 chanx_right_out[4]
rlabel metal2 24794 7837 24794 7837 0 chanx_right_out[5]
rlabel metal2 25162 8789 25162 8789 0 chanx_right_out[6]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[7]
rlabel metal2 24794 9945 24794 9945 0 chanx_right_out[8]
rlabel metal2 24794 10829 24794 10829 0 chanx_right_out[9]
rlabel metal2 1150 2438 1150 2438 0 chany_bottom_in[0]
rlabel metal2 4830 2132 4830 2132 0 chany_bottom_in[10]
rlabel metal2 5198 1894 5198 1894 0 chany_bottom_in[11]
rlabel metal2 5566 2132 5566 2132 0 chany_bottom_in[12]
rlabel metal2 5934 1894 5934 1894 0 chany_bottom_in[13]
rlabel metal2 6302 2132 6302 2132 0 chany_bottom_in[14]
rlabel metal2 6670 1588 6670 1588 0 chany_bottom_in[15]
rlabel metal2 7038 1860 7038 1860 0 chany_bottom_in[16]
rlabel metal2 7406 2132 7406 2132 0 chany_bottom_in[17]
rlabel metal2 7774 1520 7774 1520 0 chany_bottom_in[18]
rlabel metal2 8142 823 8142 823 0 chany_bottom_in[19]
rlabel metal2 1518 2098 1518 2098 0 chany_bottom_in[1]
rlabel metal2 8510 1860 8510 1860 0 chany_bottom_in[20]
rlabel metal2 8878 2438 8878 2438 0 chany_bottom_in[21]
rlabel metal2 9246 2438 9246 2438 0 chany_bottom_in[22]
rlabel metal2 9614 2132 9614 2132 0 chany_bottom_in[23]
rlabel metal2 9982 2132 9982 2132 0 chany_bottom_in[24]
rlabel metal2 10350 1860 10350 1860 0 chany_bottom_in[25]
rlabel metal2 10718 2132 10718 2132 0 chany_bottom_in[26]
rlabel metal2 11086 1792 11086 1792 0 chany_bottom_in[27]
rlabel metal2 11454 1588 11454 1588 0 chany_bottom_in[28]
rlabel metal2 11822 1860 11822 1860 0 chany_bottom_in[29]
rlabel metal2 1886 1894 1886 1894 0 chany_bottom_in[2]
rlabel metal2 2254 1588 2254 1588 0 chany_bottom_in[3]
rlabel metal2 2622 1588 2622 1588 0 chany_bottom_in[4]
rlabel metal2 2990 1299 2990 1299 0 chany_bottom_in[5]
rlabel metal2 3358 1894 3358 1894 0 chany_bottom_in[6]
rlabel metal2 3726 1894 3726 1894 0 chany_bottom_in[7]
rlabel metal2 4094 1588 4094 1588 0 chany_bottom_in[8]
rlabel metal2 4462 1894 4462 1894 0 chany_bottom_in[9]
rlabel metal2 12190 1554 12190 1554 0 chany_bottom_out[0]
rlabel metal2 15870 1860 15870 1860 0 chany_bottom_out[10]
rlabel metal2 16238 2404 16238 2404 0 chany_bottom_out[11]
rlabel metal2 16606 1826 16606 1826 0 chany_bottom_out[12]
rlabel metal2 16974 1588 16974 1588 0 chany_bottom_out[13]
rlabel metal2 17342 1792 17342 1792 0 chany_bottom_out[14]
rlabel metal2 17710 2166 17710 2166 0 chany_bottom_out[15]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out[16]
rlabel metal2 18446 823 18446 823 0 chany_bottom_out[17]
rlabel metal2 18814 1792 18814 1792 0 chany_bottom_out[18]
rlabel metal2 19182 2098 19182 2098 0 chany_bottom_out[19]
rlabel metal2 12558 2166 12558 2166 0 chany_bottom_out[1]
rlabel metal2 19550 2948 19550 2948 0 chany_bottom_out[20]
rlabel metal2 19918 1826 19918 1826 0 chany_bottom_out[21]
rlabel metal2 20286 2404 20286 2404 0 chany_bottom_out[22]
rlabel metal2 20654 3254 20654 3254 0 chany_bottom_out[23]
rlabel metal2 21022 1792 21022 1792 0 chany_bottom_out[24]
rlabel metal2 21390 1435 21390 1435 0 chany_bottom_out[25]
rlabel metal2 21758 3186 21758 3186 0 chany_bottom_out[26]
rlabel metal2 22126 1979 22126 1979 0 chany_bottom_out[27]
rlabel metal1 22540 7310 22540 7310 0 chany_bottom_out[28]
rlabel metal2 22862 2064 22862 2064 0 chany_bottom_out[29]
rlabel metal2 12926 1435 12926 1435 0 chany_bottom_out[2]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out[3]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out[4]
rlabel metal2 14030 2166 14030 2166 0 chany_bottom_out[5]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out[6]
rlabel metal2 14766 1860 14766 1860 0 chany_bottom_out[7]
rlabel metal2 15134 1622 15134 1622 0 chany_bottom_out[8]
rlabel metal2 15502 2166 15502 2166 0 chany_bottom_out[9]
rlabel metal1 12512 52462 12512 52462 0 chany_top_in_0[0]
rlabel metal1 16721 54162 16721 54162 0 chany_top_in_0[10]
rlabel metal1 16468 53550 16468 53550 0 chany_top_in_0[11]
rlabel metal1 17112 53550 17112 53550 0 chany_top_in_0[12]
rlabel metal1 17434 54230 17434 54230 0 chany_top_in_0[13]
rlabel metal1 17986 54162 17986 54162 0 chany_top_in_0[14]
rlabel metal1 17986 53550 17986 53550 0 chany_top_in_0[15]
rlabel metal2 18262 55711 18262 55711 0 chany_top_in_0[16]
rlabel metal1 19044 54162 19044 54162 0 chany_top_in_0[17]
rlabel metal1 19228 53550 19228 53550 0 chany_top_in_0[18]
rlabel metal1 19458 54230 19458 54230 0 chany_top_in_0[19]
rlabel metal1 13570 53142 13570 53142 0 chany_top_in_0[1]
rlabel metal1 19872 53074 19872 53074 0 chany_top_in_0[20]
rlabel metal1 20516 54230 20516 54230 0 chany_top_in_0[21]
rlabel metal1 20516 53550 20516 53550 0 chany_top_in_0[22]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[23]
rlabel metal1 21712 54162 21712 54162 0 chany_top_in_0[24]
rlabel metal1 21896 53550 21896 53550 0 chany_top_in_0[25]
rlabel metal1 21988 53074 21988 53074 0 chany_top_in_0[26]
rlabel metal1 22632 53074 22632 53074 0 chany_top_in_0[27]
rlabel metal2 22678 55711 22678 55711 0 chany_top_in_0[28]
rlabel metal2 23230 56236 23230 56236 0 chany_top_in_0[29]
rlabel metal2 13294 56236 13294 56236 0 chany_top_in_0[2]
rlabel metal1 13524 53074 13524 53074 0 chany_top_in_0[3]
rlabel metal1 13800 53550 13800 53550 0 chany_top_in_0[4]
rlabel metal1 14260 53550 14260 53550 0 chany_top_in_0[5]
rlabel metal1 14628 54162 14628 54162 0 chany_top_in_0[6]
rlabel metal1 15226 54230 15226 54230 0 chany_top_in_0[7]
rlabel metal1 15824 54162 15824 54162 0 chany_top_in_0[8]
rlabel metal1 15732 53550 15732 53550 0 chany_top_in_0[9]
rlabel metal2 1334 55711 1334 55711 0 chany_top_out_0[0]
rlabel metal1 5060 51918 5060 51918 0 chany_top_out_0[10]
rlabel metal1 4324 54230 4324 54230 0 chany_top_out_0[11]
rlabel metal2 5750 54682 5750 54682 0 chany_top_out_0[12]
rlabel metal2 6118 54376 6118 54376 0 chany_top_out_0[13]
rlabel metal2 6486 54342 6486 54342 0 chany_top_out_0[14]
rlabel metal2 6854 55711 6854 55711 0 chany_top_out_0[15]
rlabel metal2 6854 54281 6854 54281 0 chany_top_out_0[16]
rlabel metal1 7084 53618 7084 53618 0 chany_top_out_0[17]
rlabel metal2 7958 55711 7958 55711 0 chany_top_out_0[18]
rlabel metal2 8326 54920 8326 54920 0 chany_top_out_0[19]
rlabel metal1 1978 49742 1978 49742 0 chany_top_out_0[1]
rlabel metal2 8694 54614 8694 54614 0 chany_top_out_0[20]
rlabel metal1 9384 53618 9384 53618 0 chany_top_out_0[21]
rlabel metal1 8924 54230 8924 54230 0 chany_top_out_0[22]
rlabel metal1 10074 52530 10074 52530 0 chany_top_out_0[23]
rlabel metal1 10212 53006 10212 53006 0 chany_top_out_0[24]
rlabel metal2 10534 54920 10534 54920 0 chany_top_out_0[25]
rlabel metal2 10902 55226 10902 55226 0 chany_top_out_0[26]
rlabel metal1 11730 53006 11730 53006 0 chany_top_out_0[27]
rlabel metal1 11914 53618 11914 53618 0 chany_top_out_0[28]
rlabel metal1 12282 54094 12282 54094 0 chany_top_out_0[29]
rlabel metal1 2760 52666 2760 52666 0 chany_top_out_0[2]
rlabel metal2 2622 56236 2622 56236 0 chany_top_out_0[3]
rlabel metal2 2806 55711 2806 55711 0 chany_top_out_0[4]
rlabel metal2 3174 55711 3174 55711 0 chany_top_out_0[5]
rlabel metal2 3542 54070 3542 54070 0 chany_top_out_0[6]
rlabel metal2 4048 53244 4048 53244 0 chany_top_out_0[7]
rlabel metal1 4140 53142 4140 53142 0 chany_top_out_0[8]
rlabel metal1 3956 53618 3956 53618 0 chany_top_out_0[9]
rlabel metal1 7498 22712 7498 22712 0 clknet_0_prog_clk
rlabel metal1 5382 8602 5382 8602 0 clknet_4_0_0_prog_clk
rlabel metal1 4002 48586 4002 48586 0 clknet_4_10_0_prog_clk
rlabel metal2 11822 43214 11822 43214 0 clknet_4_11_0_prog_clk
rlabel metal1 18630 35700 18630 35700 0 clknet_4_12_0_prog_clk
rlabel metal1 20562 33966 20562 33966 0 clknet_4_13_0_prog_clk
rlabel metal1 18630 41174 18630 41174 0 clknet_4_14_0_prog_clk
rlabel metal1 23322 42228 23322 42228 0 clknet_4_15_0_prog_clk
rlabel metal2 11270 11424 11270 11424 0 clknet_4_1_0_prog_clk
rlabel metal1 2070 23732 2070 23732 0 clknet_4_2_0_prog_clk
rlabel metal1 12098 22542 12098 22542 0 clknet_4_3_0_prog_clk
rlabel metal1 17066 11730 17066 11730 0 clknet_4_4_0_prog_clk
rlabel metal1 18676 10778 18676 10778 0 clknet_4_5_0_prog_clk
rlabel metal1 14536 24786 14536 24786 0 clknet_4_6_0_prog_clk
rlabel metal1 23046 20434 23046 20434 0 clknet_4_7_0_prog_clk
rlabel metal2 7774 32912 7774 32912 0 clknet_4_8_0_prog_clk
rlabel metal1 9982 30770 9982 30770 0 clknet_4_9_0_prog_clk
rlabel metal2 2806 13617 2806 13617 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 15708 1004 15708 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18020 1004 18020 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 20332 1004 20332 0 gfpga_pad_io_soc_dir[3]
rlabel metal3 820 31892 820 31892 0 gfpga_pad_io_soc_in[0]
rlabel metal3 1234 34204 1234 34204 0 gfpga_pad_io_soc_in[1]
rlabel metal3 820 36516 820 36516 0 gfpga_pad_io_soc_in[2]
rlabel metal3 820 38828 820 38828 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 22644 1004 22644 0 gfpga_pad_io_soc_out[0]
rlabel metal3 1004 24956 1004 24956 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 27268 1004 27268 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 29580 1004 29580 0 gfpga_pad_io_soc_out[3]
rlabel metal3 1188 41140 1188 41140 0 isol_n
rlabel metal1 4140 48790 4140 48790 0 net1
rlabel metal1 19504 35054 19504 35054 0 net10
rlabel metal1 15732 17306 15732 17306 0 net100
rlabel metal1 25346 47974 25346 47974 0 net101
rlabel metal1 25208 48518 25208 48518 0 net102
rlabel metal1 19918 41242 19918 41242 0 net103
rlabel metal1 25530 50150 25530 50150 0 net104
rlabel metal1 25484 50694 25484 50694 0 net105
rlabel metal1 25438 51238 25438 51238 0 net106
rlabel metal1 24702 51782 24702 51782 0 net107
rlabel metal1 24610 5610 24610 5610 0 net108
rlabel metal1 10028 42534 10028 42534 0 net109
rlabel metal2 17710 38590 17710 38590 0 net11
rlabel metal1 2898 48042 2898 48042 0 net110
rlabel metal1 1886 50796 1886 50796 0 net111
rlabel metal2 6072 45540 6072 45540 0 net112
rlabel metal1 20102 6324 20102 6324 0 net113
rlabel metal1 4784 50286 4784 50286 0 net114
rlabel metal2 22402 12036 22402 12036 0 net115
rlabel metal1 21528 12410 21528 12410 0 net116
rlabel metal1 23920 11730 23920 11730 0 net117
rlabel metal1 22494 16626 22494 16626 0 net118
rlabel metal2 22218 16524 22218 16524 0 net119
rlabel metal1 23506 37094 23506 37094 0 net12
rlabel metal1 23736 13906 23736 13906 0 net120
rlabel metal1 21942 15504 21942 15504 0 net121
rlabel metal1 24518 18598 24518 18598 0 net122
rlabel metal1 22678 16524 22678 16524 0 net123
rlabel metal1 20286 18292 20286 18292 0 net124
rlabel metal1 24426 5202 24426 5202 0 net125
rlabel metal1 22494 17646 22494 17646 0 net126
rlabel metal1 20700 19346 20700 19346 0 net127
rlabel metal1 22402 22950 22402 22950 0 net128
rlabel metal1 24058 19822 24058 19822 0 net129
rlabel metal1 16008 37230 16008 37230 0 net13
rlabel metal1 24610 19346 24610 19346 0 net130
rlabel metal1 23552 21998 23552 21998 0 net131
rlabel metal1 23230 23086 23230 23086 0 net132
rlabel metal1 22310 23732 22310 23732 0 net133
rlabel metal1 23644 24174 23644 24174 0 net134
rlabel metal2 24150 24412 24150 24412 0 net135
rlabel metal1 23368 8806 23368 8806 0 net136
rlabel metal1 24380 8806 24380 8806 0 net137
rlabel metal1 23092 7854 23092 7854 0 net138
rlabel metal1 24380 7378 24380 7378 0 net139
rlabel metal1 17986 24242 17986 24242 0 net14
rlabel metal1 23920 8466 23920 8466 0 net140
rlabel metal1 23736 10030 23736 10030 0 net141
rlabel metal1 23782 9554 23782 9554 0 net142
rlabel metal2 23966 11084 23966 11084 0 net143
rlabel metal2 9798 8670 9798 8670 0 net144
rlabel metal1 16790 3026 16790 3026 0 net145
rlabel metal1 16054 4114 16054 4114 0 net146
rlabel metal1 18308 3026 18308 3026 0 net147
rlabel metal1 17664 2346 17664 2346 0 net148
rlabel metal2 17480 14348 17480 14348 0 net149
rlabel metal2 13018 39134 13018 39134 0 net15
rlabel metal1 18630 3502 18630 3502 0 net150
rlabel metal1 18446 12138 18446 12138 0 net151
rlabel metal1 21758 2414 21758 2414 0 net152
rlabel metal1 19412 4590 19412 4590 0 net153
rlabel metal1 20930 7786 20930 7786 0 net154
rlabel metal1 12466 3468 12466 3468 0 net155
rlabel metal2 19642 8636 19642 8636 0 net156
rlabel metal1 20930 4590 20930 4590 0 net157
rlabel metal1 21850 4182 21850 4182 0 net158
rlabel metal1 19734 8874 19734 8874 0 net159
rlabel metal1 19918 32198 19918 32198 0 net16
rlabel metal1 19090 6698 19090 6698 0 net160
rlabel metal1 23322 5542 23322 5542 0 net161
rlabel metal1 21528 5814 21528 5814 0 net162
rlabel metal1 21068 5882 21068 5882 0 net163
rlabel metal1 20240 6426 20240 6426 0 net164
rlabel metal1 20148 6630 20148 6630 0 net165
rlabel metal1 13432 4114 13432 4114 0 net166
rlabel metal1 12052 2482 12052 2482 0 net167
rlabel metal1 12742 3026 12742 3026 0 net168
rlabel metal1 14076 12682 14076 12682 0 net169
rlabel metal1 19550 34646 19550 34646 0 net17
rlabel metal1 15502 2414 15502 2414 0 net170
rlabel metal2 14858 6460 14858 6460 0 net171
rlabel metal1 16836 2414 16836 2414 0 net172
rlabel metal1 15640 13226 15640 13226 0 net173
rlabel metal2 1610 44948 1610 44948 0 net174
rlabel metal1 5566 51986 5566 51986 0 net175
rlabel metal1 5336 51578 5336 51578 0 net176
rlabel metal1 5612 53074 5612 53074 0 net177
rlabel metal1 5612 52462 5612 52462 0 net178
rlabel metal1 7958 43962 7958 43962 0 net179
rlabel metal1 23736 41582 23736 41582 0 net18
rlabel metal2 7130 51238 7130 51238 0 net180
rlabel metal1 5865 54162 5865 54162 0 net181
rlabel metal2 5382 44105 5382 44105 0 net182
rlabel metal1 9430 43962 9430 43962 0 net183
rlabel metal1 7636 49946 7636 49946 0 net184
rlabel metal1 2852 42330 2852 42330 0 net185
rlabel metal1 9982 43894 9982 43894 0 net186
rlabel metal1 9660 45050 9660 45050 0 net187
rlabel metal1 9752 45390 9752 45390 0 net188
rlabel metal2 9614 51170 9614 51170 0 net189
rlabel metal1 25208 42534 25208 42534 0 net19
rlabel metal2 9430 51748 9430 51748 0 net190
rlabel metal1 10442 44302 10442 44302 0 net191
rlabel metal2 9890 52598 9890 52598 0 net192
rlabel metal2 10534 52054 10534 52054 0 net193
rlabel metal2 11730 52836 11730 52836 0 net194
rlabel metal1 11960 52666 11960 52666 0 net195
rlabel metal1 2898 50286 2898 50286 0 net196
rlabel metal1 2254 51306 2254 51306 0 net197
rlabel metal1 4094 42738 4094 42738 0 net198
rlabel metal1 4002 41786 4002 41786 0 net199
rlabel metal1 2576 3706 2576 3706 0 net2
rlabel metal1 25346 43622 25346 43622 0 net20
rlabel metal1 5612 41718 5612 41718 0 net200
rlabel metal1 4186 51374 4186 51374 0 net201
rlabel metal1 6532 42738 6532 42738 0 net202
rlabel metal2 6578 44751 6578 44751 0 net203
rlabel metal1 2208 13906 2208 13906 0 net204
rlabel metal1 1932 18598 1932 18598 0 net205
rlabel metal1 1840 18258 1840 18258 0 net206
rlabel metal2 1794 21148 1794 21148 0 net207
rlabel metal2 2714 22644 2714 22644 0 net208
rlabel metal1 1886 22746 1886 22746 0 net209
rlabel metal1 24288 43214 24288 43214 0 net21
rlabel metal1 2024 24650 2024 24650 0 net210
rlabel metal1 1932 27098 1932 27098 0 net211
rlabel metal1 17986 5202 17986 5202 0 net212
rlabel metal2 24610 45254 24610 45254 0 net213
rlabel metal2 23782 53380 23782 53380 0 net214
rlabel metal1 22310 8500 22310 8500 0 net215
rlabel metal1 25070 53074 25070 53074 0 net216
rlabel metal1 22816 6086 22816 6086 0 net217
rlabel metal1 22862 53516 22862 53516 0 net218
rlabel metal1 17112 20570 17112 20570 0 net219
rlabel metal2 24978 42942 24978 42942 0 net22
rlabel metal1 13156 27438 13156 27438 0 net220
rlabel metal1 23276 31926 23276 31926 0 net221
rlabel metal1 23046 20910 23046 20910 0 net222
rlabel metal1 15272 36754 15272 36754 0 net223
rlabel metal1 17434 21522 17434 21522 0 net224
rlabel metal2 22218 28730 22218 28730 0 net225
rlabel metal2 16330 36346 16330 36346 0 net226
rlabel metal2 19642 37434 19642 37434 0 net227
rlabel metal1 16238 37842 16238 37842 0 net228
rlabel metal2 14030 39440 14030 39440 0 net229
rlabel metal1 18078 40358 18078 40358 0 net23
rlabel metal1 13800 37842 13800 37842 0 net230
rlabel metal2 24978 39950 24978 39950 0 net231
rlabel metal1 13386 32402 13386 32402 0 net232
rlabel metal2 10994 29818 10994 29818 0 net233
rlabel metal1 13064 25262 13064 25262 0 net234
rlabel metal2 10534 26894 10534 26894 0 net235
rlabel metal1 8418 26010 8418 26010 0 net236
rlabel metal2 9338 26758 9338 26758 0 net237
rlabel metal2 8234 24378 8234 24378 0 net238
rlabel metal1 10580 23698 10580 23698 0 net239
rlabel metal1 23782 45798 23782 45798 0 net24
rlabel metal1 6486 9554 6486 9554 0 net240
rlabel metal1 15502 11730 15502 11730 0 net241
rlabel metal1 20470 34408 20470 34408 0 net242
rlabel metal2 17250 13124 17250 13124 0 net243
rlabel metal1 18676 14994 18676 14994 0 net244
rlabel metal1 20838 15470 20838 15470 0 net245
rlabel metal2 24426 15640 24426 15640 0 net246
rlabel metal1 19596 15130 19596 15130 0 net247
rlabel metal2 23322 13736 23322 13736 0 net248
rlabel metal1 20332 11118 20332 11118 0 net249
rlabel metal1 15686 26010 15686 26010 0 net25
rlabel metal1 18676 13294 18676 13294 0 net250
rlabel metal1 23322 34578 23322 34578 0 net251
rlabel metal1 21298 40154 21298 40154 0 net252
rlabel metal1 10856 37978 10856 37978 0 net253
rlabel metal1 7912 30906 7912 30906 0 net254
rlabel metal2 8694 32572 8694 32572 0 net255
rlabel metal1 12696 38930 12696 38930 0 net256
rlabel metal1 8142 31314 8142 31314 0 net257
rlabel metal1 4830 31450 4830 31450 0 net258
rlabel metal1 8464 38318 8464 38318 0 net259
rlabel metal1 17848 25806 17848 25806 0 net26
rlabel metal2 9982 35802 9982 35802 0 net260
rlabel metal1 11500 37842 11500 37842 0 net261
rlabel metal2 15226 35598 15226 35598 0 net262
rlabel metal1 7544 30702 7544 30702 0 net263
rlabel metal2 25346 4879 25346 4879 0 net264
rlabel metal1 10396 23086 10396 23086 0 net265
rlabel metal1 11454 19822 11454 19822 0 net266
rlabel metal1 8878 16218 8878 16218 0 net267
rlabel metal1 8970 23834 8970 23834 0 net268
rlabel metal2 13754 21318 13754 21318 0 net269
rlabel metal1 19504 33354 19504 33354 0 net27
rlabel metal2 13478 24004 13478 24004 0 net270
rlabel metal2 19550 25296 19550 25296 0 net271
rlabel metal1 22356 24378 22356 24378 0 net272
rlabel metal1 17848 28526 17848 28526 0 net273
rlabel metal1 18722 34918 18722 34918 0 net28
rlabel metal1 18906 33966 18906 33966 0 net29
rlabel metal1 21206 26010 21206 26010 0 net3
rlabel metal1 22724 32538 22724 32538 0 net30
rlabel metal1 16652 36754 16652 36754 0 net31
rlabel metal1 17250 32266 17250 32266 0 net32
rlabel metal1 3588 3978 3588 3978 0 net33
rlabel metal2 5106 3944 5106 3944 0 net34
rlabel metal2 5198 4692 5198 4692 0 net35
rlabel metal2 16054 4420 16054 4420 0 net36
rlabel metal1 6072 3094 6072 3094 0 net37
rlabel metal1 6670 3706 6670 3706 0 net38
rlabel metal1 6210 2618 6210 2618 0 net39
rlabel metal1 14398 31892 14398 31892 0 net4
rlabel metal1 11224 3094 11224 3094 0 net40
rlabel metal2 7682 3927 7682 3927 0 net41
rlabel metal1 8004 2550 8004 2550 0 net42
rlabel via2 8418 3723 8418 3723 0 net43
rlabel metal1 3450 3638 3450 3638 0 net44
rlabel metal1 11040 4998 11040 4998 0 net45
rlabel metal1 7958 3978 7958 3978 0 net46
rlabel metal1 10488 44778 10488 44778 0 net47
rlabel metal1 9568 3706 9568 3706 0 net48
rlabel metal1 12558 3366 12558 3366 0 net49
rlabel metal1 23736 32742 23736 32742 0 net5
rlabel metal1 13248 5610 13248 5610 0 net50
rlabel metal2 11546 3944 11546 3944 0 net51
rlabel metal1 12834 2550 12834 2550 0 net52
rlabel metal1 13524 2618 13524 2618 0 net53
rlabel metal2 12006 4963 12006 4963 0 net54
rlabel metal2 2162 4352 2162 4352 0 net55
rlabel metal2 2070 4148 2070 4148 0 net56
rlabel metal1 2622 2312 2622 2312 0 net57
rlabel metal1 3358 3706 3358 3706 0 net58
rlabel metal1 3496 3094 3496 3094 0 net59
rlabel metal2 20838 30804 20838 30804 0 net6
rlabel metal1 5520 2890 5520 2890 0 net60
rlabel metal1 5681 2482 5681 2482 0 net61
rlabel metal2 5106 2873 5106 2873 0 net62
rlabel metal1 12972 52598 12972 52598 0 net63
rlabel metal1 16422 54026 16422 54026 0 net64
rlabel metal1 16468 53414 16468 53414 0 net65
rlabel metal2 17250 50048 17250 50048 0 net66
rlabel via3 17365 20604 17365 20604 0 net67
rlabel metal3 17963 20468 17963 20468 0 net68
rlabel metal1 18354 53482 18354 53482 0 net69
rlabel metal1 19412 32538 19412 32538 0 net7
rlabel metal1 18630 46682 18630 46682 0 net70
rlabel metal1 18216 12070 18216 12070 0 net71
rlabel metal1 19872 53414 19872 53414 0 net72
rlabel metal1 20562 54026 20562 54026 0 net73
rlabel via3 14605 52564 14605 52564 0 net74
rlabel metal1 19872 46002 19872 46002 0 net75
rlabel metal1 19504 12138 19504 12138 0 net76
rlabel metal1 21574 53448 21574 53448 0 net77
rlabel metal1 19872 13974 19872 13974 0 net78
rlabel metal1 21942 53958 21942 53958 0 net79
rlabel metal1 20194 36312 20194 36312 0 net8
rlabel metal1 21666 45934 21666 45934 0 net80
rlabel metal3 22287 52564 22287 52564 0 net81
rlabel metal2 22770 47226 22770 47226 0 net82
rlabel metal1 22770 44778 22770 44778 0 net83
rlabel metal1 23966 53414 23966 53414 0 net84
rlabel metal1 13800 52462 13800 52462 0 net85
rlabel metal1 10350 23528 10350 23528 0 net86
rlabel metal1 13064 53414 13064 53414 0 net87
rlabel metal1 13478 12138 13478 12138 0 net88
rlabel metal1 10718 22950 10718 22950 0 net89
rlabel metal1 23138 32878 23138 32878 0 net9
rlabel metal3 15847 21692 15847 21692 0 net90
rlabel metal1 17710 47056 17710 47056 0 net91
rlabel metal1 15410 12138 15410 12138 0 net92
rlabel metal1 2806 26418 2806 26418 0 net93
rlabel metal1 3680 27506 3680 27506 0 net94
rlabel metal1 3726 28594 3726 28594 0 net95
rlabel metal1 1748 38726 1748 38726 0 net96
rlabel metal2 4002 24922 4002 24922 0 net97
rlabel metal1 4278 23766 4278 23766 0 net98
rlabel metal1 24104 6698 24104 6698 0 net99
rlabel metal2 23230 1639 23230 1639 0 prog_clk
rlabel metal2 23598 1894 23598 1894 0 prog_reset_bottom_in
rlabel metal2 23966 1928 23966 1928 0 prog_reset_bottom_out
rlabel metal3 25584 45764 25584 45764 0 prog_reset_right_out
rlabel metal1 24012 54230 24012 54230 0 prog_reset_top_out
rlabel metal2 24334 2098 24334 2098 0 reset_bottom_in
rlabel metal2 24702 2115 24702 2115 0 reset_bottom_out
rlabel metal2 24886 54682 24886 54682 0 reset_top_out
rlabel metal2 25070 47379 25070 47379 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 25070 47957 25070 47957 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 25070 48603 25070 48603 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel via2 25070 49181 25070 49181 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25070 50065 25070 50065 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 25070 50711 25070 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 25070 51289 25070 51289 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 25162 51935 25162 51935 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1970 4148 1970 4148 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1924 6460 1924 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1878 8772 1878 8772 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1740 11084 1740 11084 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18676 14042 18676 14042 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal2 16054 20570 16054 20570 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 12558 21012 12558 21012 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 15410 22746 15410 22746 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 18814 21012 18814 21012 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal2 16330 24956 16330 24956 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 18630 32266 18630 32266 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 16514 26554 16514 26554 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 20930 24684 20930 24684 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 17986 29682 17986 29682 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20608 26894 20608 26894 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal2 22494 25908 22494 25908 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 20332 26418 20332 26418 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal1 23920 27574 23920 27574 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 15870 28730 15870 28730 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 19320 33014 19320 33014 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 16192 28594 16192 28594 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal1 20654 20230 20654 20230 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 18400 26894 18400 26894 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 18584 22746 18584 22746 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 16698 32810 16698 32810 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 15778 32334 15778 32334 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 15410 32198 15410 32198 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal2 21022 33626 21022 33626 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 20792 34034 20792 34034 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal2 23138 32895 23138 32895 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 22586 20298 22586 20298 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal2 21298 23392 21298 23392 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 23690 20536 23690 20536 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 12282 43112 12282 43112 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 23828 21454 23828 21454 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal2 19918 21726 19918 21726 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 18860 35734 18860 35734 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 24472 30022 24472 30022 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal1 21160 31858 21160 31858 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 22586 30124 22586 30124 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 23138 43622 23138 43622 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 20148 40902 20148 40902 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 20286 39474 20286 39474 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal2 18722 38658 18722 38658 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 19596 42330 19596 42330 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal1 19780 44778 19780 44778 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 20010 40528 20010 40528 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 17802 39474 17802 39474 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 18722 45492 18722 45492 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal2 16330 39893 16330 39893 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal2 16054 45764 16054 45764 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal2 17434 46852 17434 46852 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 14444 38862 14444 38862 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal2 16054 40131 16054 40131 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 15916 46682 15916 46682 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal2 13892 40732 13892 40732 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal2 23598 42398 23598 42398 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal2 20654 36380 20654 36380 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 25024 40902 25024 40902 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 13984 34918 13984 34918 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal1 13800 41174 13800 41174 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 15226 37774 15226 37774 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 13570 29614 13570 29614 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13202 35802 13202 35802 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal2 11270 30294 11270 30294 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal2 13570 24990 13570 24990 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal2 12834 26860 12834 26860 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal1 11040 28186 11040 28186 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 14720 30090 14720 30090 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 8188 28390 8188 28390 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal1 7498 25874 7498 25874 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 9476 25806 9476 25806 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 9016 28186 9016 28186 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 9614 24718 9614 24718 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal2 7498 24786 7498 24786 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal2 10902 23290 10902 23290 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal2 9430 24446 9430 24446 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal1 9660 12750 9660 12750 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 11684 24718 11684 24718 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 8050 17068 8050 17068 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 12926 11832 12926 11832 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 11362 11050 11362 11050 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal1 22816 36822 22816 36822 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 23782 41990 23782 41990 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal2 21666 35870 21666 35870 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 15686 12954 15686 12954 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal1 14490 11866 14490 11866 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal1 18538 16218 18538 16218 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 17158 16558 17158 16558 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 20010 17374 20010 17374 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal1 19504 17714 19504 17714 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 22954 16966 22954 16966 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 22310 17272 22310 17272 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal1 22448 16150 22448 16150 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 22494 18632 22494 18632 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 21298 13804 21298 13804 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal1 22931 15878 22931 15878 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 20010 11424 20010 11424 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal1 18952 12750 18952 12750 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 18078 11866 18078 11866 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24794 37978 24794 37978 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 20102 33456 20102 33456 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal1 23368 35122 23368 35122 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 22494 43214 22494 43214 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 22402 42126 22402 42126 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 12374 44506 12374 44506 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 10074 42772 10074 42772 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 11730 44166 11730 44166 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 6762 38522 6762 38522 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal1 6532 35802 6532 35802 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal2 7590 30498 7590 30498 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal2 10350 35326 10350 35326 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal2 9522 35122 9522 35122 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal1 9706 28628 9706 28628 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 12834 33388 12834 33388 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 11730 42058 11730 42058 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 13018 34034 13018 34034 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14398 39474 14398 39474 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal2 6946 33558 6946 33558 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal2 8050 29920 8050 29920 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 8970 30158 8970 30158 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 5750 36652 5750 36652 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 12742 34612 12742 34612 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 5290 31246 5290 31246 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal2 8510 41888 8510 41888 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 13202 39542 13202 39542 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 12558 38352 12558 38352 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal2 9338 37876 9338 37876 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 14950 38352 14950 38352 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal2 13478 36074 13478 36074 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13110 41480 13110 41480 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal1 11546 41514 11546 41514 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 17986 39032 17986 39032 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 16974 37910 16974 37910 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 8326 30770 8326 30770 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal2 7866 37264 7866 37264 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 19642 6800 19642 6800 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal2 15594 26316 15594 26316 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16100 25126 16100 25126 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11960 21114 11960 21114 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14996 20570 14996 20570 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14306 20570 14306 20570 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14766 18734 14766 18734 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 17158 6766 17158 6766 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal2 17342 29104 17342 29104 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18768 32198 18768 32198 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 24242 15870 24242 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13110 23970 13110 23970 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16376 23086 16376 23086 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15778 23086 15778 23086 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16100 16558 16100 16558 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18676 8942 18676 8942 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 19596 27982 19596 27982 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 28118 20194 28118 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 24786 19550 24786 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19918 26044 19918 26044 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 24378 19826 24378 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 18722 20713 18722 20713 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 20608 7854 20608 7854 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 19366 30090 19366 30090 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22494 28186 22494 28186 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22494 24718 22494 24718 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 25500 21942 25500 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22126 23834 22126 23834 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21114 14994 21114 14994 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16054 8942 16054 8942 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal2 17802 32028 17802 32028 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19366 34986 19366 34986 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17756 28186 17756 28186 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17296 31926 17296 31926 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17066 27438 17066 27438 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16422 20434 16422 20434 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 18400 6290 18400 6290 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal1 17940 24718 17940 24718 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18860 24922 18860 24922 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18216 24582 18216 24582 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18308 19686 18308 19686 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18078 14382 18078 14382 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14260 9622 14260 9622 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal2 16146 34782 16146 34782 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16330 32878 16330 32878 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 32742 15226 32742 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13708 27370 13708 27370 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13662 21998 13662 21998 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18584 10030 18584 10030 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 21022 36142 21022 36142 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21620 34714 21620 34714 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22448 32198 22448 32198 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20976 21692 20976 21692 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 20194 6289 20194 6289 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 21942 28424 21942 28424 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22011 29750 22011 29750 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20608 21556 20608 21556 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22540 20502 22540 20502 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22678 20570 22678 20570 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 20654 17340 20654 17340 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10212 25126 10212 25126 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 13432 37094 13432 37094 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15318 37026 15318 37026 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10948 25262 10948 25262 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16606 9605 16606 9605 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal2 19550 26792 19550 26792 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19964 25874 19964 25874 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18216 22066 18216 22066 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17894 21998 17894 21998 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 18676 22542 18676 22542 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18216 20910 18216 20910 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 16606 19754 16606 19754 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 24380 25262 24380 25262 0 sb_0__1_.mux_right_track_0.out
rlabel metal1 21206 31926 21206 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22080 31926 22080 31926 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23552 29682 23552 29682 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 29104 23322 29104 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24104 28050 24104 28050 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24104 32198 24104 32198 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 19826 41650 19826 41650 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 41446 19688 41446 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19642 38386 19642 38386 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17296 36346 17296 36346 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24058 32436 24058 32436 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 25254 28560 25254 28560 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19780 40562 19780 40562 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 39066 20056 39066 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16560 37094 16560 37094 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 19504 35292 19504 35292 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22034 29104 22034 29104 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 17940 42738 17940 42738 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17986 39406 17986 39406 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15778 38216 15778 38216 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17434 35938 17434 35938 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20562 32742 20562 32742 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 17296 43418 17296 43418 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16514 40494 16514 40494 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14950 38794 14950 38794 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 32878 19458 32878 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19964 31926 19964 31926 0 sb_0__1_.mux_right_track_18.out
rlabel metal2 17342 44064 17342 44064 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 39066 16422 39066 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14398 37978 14398 37978 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18400 31790 18400 31790 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 29206 24656 29206 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 22678 41242 22678 41242 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22126 39780 22126 39780 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20010 36210 20010 36210 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23736 40494 23736 40494 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24150 39610 24150 39610 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24794 34000 24794 34000 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 22126 27047 22126 27047 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 14812 37910 14812 37910 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15042 33626 15042 33626 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13984 33082 13984 33082 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14904 33286 14904 33286 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21068 20502 21068 20502 0 sb_0__1_.mux_right_track_22.out
rlabel metal2 13938 36295 13938 36295 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13478 31484 13478 31484 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12282 29580 12282 29580 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19642 25296 19642 25296 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 18734 24656 18734 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 14720 24242 14720 24242 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14628 24038 14628 24038 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19550 20910 19550 20910 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19688 19754 19688 19754 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 13386 26350 13386 26350 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11638 26418 11638 26418 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18354 23052 18354 23052 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16652 19482 16652 19482 0 sb_0__1_.mux_right_track_28.out
rlabel metal2 10442 28424 10442 28424 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8464 25738 8464 25738 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12052 24412 12052 24412 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22218 21182 22218 21182 0 sb_0__1_.mux_right_track_30.out
rlabel metal1 10350 26010 10350 26010 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9476 25942 9476 25942 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15318 21522 15318 21522 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21942 18258 21942 18258 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 11454 27914 11454 27914 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8694 24378 8694 24378 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14996 20978 14996 20978 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21160 16150 21160 16150 0 sb_0__1_.mux_right_track_34.out
rlabel metal2 12374 25840 12374 25840 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10994 23834 10994 23834 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16698 19346 16698 19346 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18837 12206 18837 12206 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 10810 24786 10810 24786 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9384 12954 9384 12954 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7958 12818 7958 12818 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15088 12206 15088 12206 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20378 11322 20378 11322 0 sb_0__1_.mux_right_track_38.out
rlabel metal2 14766 12240 14766 12240 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17457 11118 17457 11118 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24288 27438 24288 27438 0 sb_0__1_.mux_right_track_4.out
rlabel metal2 21666 42092 21666 42092 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22310 38896 22310 38896 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22632 35666 22632 35666 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19090 34476 19090 34476 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 22770 33677 22770 33677 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 11764 23414 11764 0 sb_0__1_.mux_right_track_40.out
rlabel metal2 17342 13498 17342 13498 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 11730 19688 11730 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 12206 24702 12206 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 18216 15470 18216 15470 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22264 13906 22264 13906 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 11152 24058 11152 0 sb_0__1_.mux_right_track_46.out
rlabel metal2 20470 17544 20470 17544 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 13872 22862 13872 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24794 10064 24794 10064 0 sb_0__1_.mux_right_track_48.out
rlabel metal1 21068 15334 21068 15334 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23966 14450 23966 14450 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24058 11050 24058 11050 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21620 18734 21620 18734 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19182 15130 19182 15130 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22310 18258 22310 18258 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24794 8976 24794 8976 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 21114 14042 21114 14042 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22402 11118 22402 11118 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24058 9146 24058 9146 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 19826 11186 19826 11186 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 10404 22218 10404 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24794 7854 24794 7854 0 sb_0__1_.mux_right_track_56.out
rlabel metal1 18492 13362 18492 13362 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19734 13498 19734 13498 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 31926 24656 31926 0 sb_0__1_.mux_right_track_6.out
rlabel metal2 21574 39882 21574 39882 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21482 37298 21482 37298 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 33626 20148 33626 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23736 36210 23736 36210 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23276 35258 23276 35258 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24794 31824 24794 31824 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24196 28118 24196 28118 0 sb_0__1_.mux_right_track_8.out
rlabel metal2 22494 44200 22494 44200 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20746 40902 20746 40902 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 37094 19688 37094 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21988 41990 21988 41990 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20746 40120 20746 40120 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 23874 37060 23874 37060 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11868 48858 11868 48858 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 9430 42568 9430 42568 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 40698 16284 40698 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15180 35802 15180 35802 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11132 37706 11132 37706 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12236 43418 12236 43418 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12052 44370 12052 44370 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11822 48722 11822 48722 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7406 44234 7406 44234 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 9522 37230 9522 37230 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16882 36312 16882 36312 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11546 30090 11546 30090 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8188 33626 8188 33626 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9016 37094 9016 37094 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9936 33626 9936 33626 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7912 44370 7912 44370 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8510 42534 8510 42534 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 12788 33626 12788 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16054 33558 16054 33558 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9246 28730 9246 28730 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11270 33626 11270 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9246 33082 9246 33082 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7406 42602 7406 42602 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11730 47226 11730 47226 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 14996 39406 14996 39406 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18584 35190 18584 35190 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12098 34170 12098 34170 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12236 42262 12236 42262 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12006 42194 12006 42194 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11684 42330 11684 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 7038 44037 7038 44037 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 12144 32742 12144 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15134 29750 15134 29750 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9062 29818 9062 29818 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10672 33082 10672 33082 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 7682 31994 7682 31994 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7176 42670 7176 42670 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 5980 50286 5980 50286 0 sb_0__1_.mux_top_track_28.out
rlabel metal2 12466 34986 12466 34986 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12190 31994 12190 31994 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9154 35530 9154 35530 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 4600 31450 4600 31450 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5474 43282 5474 43282 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 6118 51340 6118 51340 0 sb_0__1_.mux_top_track_36.out
rlabel metal2 12374 38828 12374 38828 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8970 41446 8970 41446 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8050 41446 8050 41446 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7544 46546 7544 46546 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9890 45322 9890 45322 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 13892 36890 13892 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16376 33354 16376 33354 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10120 31450 10120 31450 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12834 36890 12834 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9844 35258 9844 35258 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10028 44166 10028 44166 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 6854 50150 6854 50150 0 sb_0__1_.mux_top_track_44.out
rlabel metal1 16376 42602 16376 42602 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11960 42602 11960 42602 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11316 42534 11316 42534 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9108 45526 9108 45526 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 21114 36890 21114 36890 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19504 36890 19504 36890 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 35258 15226 35258 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11178 45492 11178 45492 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9108 50898 9108 50898 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 9890 38250 9890 38250 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16974 36278 16974 36278 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12650 30838 12650 30838 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7406 30838 7406 30838 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9476 38522 9476 38522 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8372 34714 8372 34714 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8142 45458 8142 45458 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 25070 1826 25070 1826 0 test_enable_bottom_in
rlabel metal1 23368 7446 23368 7446 0 test_enable_bottom_out
rlabel metal1 24748 53618 24748 53618 0 test_enable_top_out
rlabel metal3 820 45764 820 45764 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 820 48076 820 48076 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 820 50388 820 50388 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1004 52700 1004 52700 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
