magic
tech sky130A
magscale 1 2
timestamp 1656241649
<< obsli1 >>
rect 1104 2159 23460 22321
<< obsm1 >>
rect 290 2128 24182 22840
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 15106 23800 15162 24600
rect 15750 23800 15806 24600
rect 16394 23800 16450 24600
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21546 23800 21602 24600
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 2134 0 2190 800
rect 6182 0 6238 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18326 0 18382 800
rect 22374 0 22430 800
<< obsm2 >>
rect 406 23744 882 23882
rect 1050 23744 1526 23882
rect 1694 23744 2170 23882
rect 2338 23744 2814 23882
rect 2982 23744 3458 23882
rect 3626 23744 4102 23882
rect 4270 23744 4746 23882
rect 4914 23744 5390 23882
rect 5558 23744 6034 23882
rect 6202 23744 6678 23882
rect 6846 23744 7322 23882
rect 7490 23744 7966 23882
rect 8134 23744 8610 23882
rect 8778 23744 9254 23882
rect 9422 23744 9898 23882
rect 10066 23744 10542 23882
rect 10710 23744 11186 23882
rect 11354 23744 11830 23882
rect 11998 23744 12474 23882
rect 12642 23744 13118 23882
rect 13286 23744 13762 23882
rect 13930 23744 14406 23882
rect 14574 23744 15050 23882
rect 15218 23744 15694 23882
rect 15862 23744 16338 23882
rect 16506 23744 16982 23882
rect 17150 23744 17626 23882
rect 17794 23744 18270 23882
rect 18438 23744 18914 23882
rect 19082 23744 19558 23882
rect 19726 23744 20202 23882
rect 20370 23744 20846 23882
rect 21014 23744 21490 23882
rect 21658 23744 22134 23882
rect 22302 23744 22778 23882
rect 22946 23744 23422 23882
rect 23590 23744 24066 23882
rect 296 856 24176 23744
rect 296 800 2078 856
rect 2246 800 6126 856
rect 6294 800 10174 856
rect 10342 800 14222 856
rect 14390 800 18270 856
rect 18438 800 22318 856
rect 22486 800 24176 856
<< metal3 >>
rect 23800 22040 24600 22160
rect 0 21360 800 21480
rect 23800 21496 24600 21616
rect 23800 20952 24600 21072
rect 23800 20408 24600 20528
rect 23800 19864 24600 19984
rect 23800 19320 24600 19440
rect 23800 18776 24600 18896
rect 23800 18232 24600 18352
rect 23800 17688 24600 17808
rect 23800 17144 24600 17264
rect 23800 16600 24600 16720
rect 23800 16056 24600 16176
rect 23800 15512 24600 15632
rect 0 15240 800 15360
rect 23800 14968 24600 15088
rect 23800 14424 24600 14544
rect 23800 13880 24600 14000
rect 23800 13336 24600 13456
rect 23800 12792 24600 12912
rect 23800 12248 24600 12368
rect 23800 11704 24600 11824
rect 23800 11160 24600 11280
rect 23800 10616 24600 10736
rect 23800 10072 24600 10192
rect 23800 9528 24600 9648
rect 0 9120 800 9240
rect 23800 8984 24600 9104
rect 23800 8440 24600 8560
rect 23800 7896 24600 8016
rect 23800 7352 24600 7472
rect 23800 6808 24600 6928
rect 23800 6264 24600 6384
rect 23800 5720 24600 5840
rect 23800 5176 24600 5296
rect 23800 4632 24600 4752
rect 23800 4088 24600 4208
rect 23800 3544 24600 3664
rect 0 3000 800 3120
rect 23800 3000 24600 3120
rect 23800 2456 24600 2576
<< obsm3 >>
rect 800 22240 23800 22337
rect 800 21960 23720 22240
rect 800 21696 23800 21960
rect 800 21560 23720 21696
rect 880 21416 23720 21560
rect 880 21280 23800 21416
rect 800 21152 23800 21280
rect 800 20872 23720 21152
rect 800 20608 23800 20872
rect 800 20328 23720 20608
rect 800 20064 23800 20328
rect 800 19784 23720 20064
rect 800 19520 23800 19784
rect 800 19240 23720 19520
rect 800 18976 23800 19240
rect 800 18696 23720 18976
rect 800 18432 23800 18696
rect 800 18152 23720 18432
rect 800 17888 23800 18152
rect 800 17608 23720 17888
rect 800 17344 23800 17608
rect 800 17064 23720 17344
rect 800 16800 23800 17064
rect 800 16520 23720 16800
rect 800 16256 23800 16520
rect 800 15976 23720 16256
rect 800 15712 23800 15976
rect 800 15440 23720 15712
rect 880 15432 23720 15440
rect 880 15168 23800 15432
rect 880 15160 23720 15168
rect 800 14888 23720 15160
rect 800 14624 23800 14888
rect 800 14344 23720 14624
rect 800 14080 23800 14344
rect 800 13800 23720 14080
rect 800 13536 23800 13800
rect 800 13256 23720 13536
rect 800 12992 23800 13256
rect 800 12712 23720 12992
rect 800 12448 23800 12712
rect 800 12168 23720 12448
rect 800 11904 23800 12168
rect 800 11624 23720 11904
rect 800 11360 23800 11624
rect 800 11080 23720 11360
rect 800 10816 23800 11080
rect 800 10536 23720 10816
rect 800 10272 23800 10536
rect 800 9992 23720 10272
rect 800 9728 23800 9992
rect 800 9448 23720 9728
rect 800 9320 23800 9448
rect 880 9184 23800 9320
rect 880 9040 23720 9184
rect 800 8904 23720 9040
rect 800 8640 23800 8904
rect 800 8360 23720 8640
rect 800 8096 23800 8360
rect 800 7816 23720 8096
rect 800 7552 23800 7816
rect 800 7272 23720 7552
rect 800 7008 23800 7272
rect 800 6728 23720 7008
rect 800 6464 23800 6728
rect 800 6184 23720 6464
rect 800 5920 23800 6184
rect 800 5640 23720 5920
rect 800 5376 23800 5640
rect 800 5096 23720 5376
rect 800 4832 23800 5096
rect 800 4552 23720 4832
rect 800 4288 23800 4552
rect 800 4008 23720 4288
rect 800 3744 23800 4008
rect 800 3464 23720 3744
rect 800 3200 23800 3464
rect 880 2920 23720 3200
rect 800 2656 23800 2920
rect 800 2376 23720 2656
rect 800 2143 23800 2376
<< metal4 >>
rect 3743 2128 4063 22352
rect 6542 2128 6862 22352
rect 9341 2128 9661 22352
rect 12140 2128 12460 22352
rect 14939 2128 15259 22352
rect 17738 2128 18058 22352
rect 20537 2128 20857 22352
<< obsm4 >>
rect 13859 4387 14859 22133
rect 15339 4387 17658 22133
rect 18138 4387 20457 22133
rect 20937 4387 21653 22133
<< labels >>
rlabel metal2 s 17038 23800 17094 24600 6 SC_IN_TOP
port 1 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 SC_OUT_BOT
port 2 nsew signal output
rlabel metal2 s 17682 23800 17738 24600 6 SC_OUT_TOP
port 3 nsew signal output
rlabel metal3 s 23800 7896 24600 8016 6 Test_en_E_in
port 4 nsew signal input
rlabel metal3 s 23800 7352 24600 7472 6 Test_en_E_out
port 5 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 Test_en_W_in
port 6 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 Test_en_W_out
port 7 nsew signal output
rlabel metal4 s 6542 2128 6862 22352 6 VGND
port 8 nsew ground bidirectional
rlabel metal4 s 12140 2128 12460 22352 6 VGND
port 8 nsew ground bidirectional
rlabel metal4 s 17738 2128 18058 22352 6 VGND
port 8 nsew ground bidirectional
rlabel metal4 s 3743 2128 4063 22352 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 9341 2128 9661 22352 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 14939 2128 15259 22352 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 20537 2128 20857 22352 6 VPWR
port 9 nsew power bidirectional
rlabel metal2 s 2134 0 2190 800 6 bottom_width_0_height_0__pin_50_
port 10 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 bottom_width_0_height_0__pin_51_
port 11 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 ccff_head
port 12 nsew signal input
rlabel metal3 s 23800 6808 24600 6928 6 ccff_tail
port 13 nsew signal output
rlabel metal2 s 18326 23800 18382 24600 6 clk_0_N_in
port 14 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 clk_0_S_in
port 15 nsew signal input
rlabel metal3 s 23800 8984 24600 9104 6 prog_clk_0_E_out
port 16 nsew signal output
rlabel metal3 s 23800 8440 24600 8560 6 prog_clk_0_N_in
port 17 nsew signal input
rlabel metal2 s 18970 23800 19026 24600 6 prog_clk_0_N_out
port 18 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 prog_clk_0_S_in
port 19 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 prog_clk_0_S_out
port 20 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 prog_clk_0_W_out
port 21 nsew signal output
rlabel metal3 s 23800 9528 24600 9648 6 right_width_0_height_0__pin_16_
port 22 nsew signal input
rlabel metal3 s 23800 10072 24600 10192 6 right_width_0_height_0__pin_17_
port 23 nsew signal input
rlabel metal3 s 23800 10616 24600 10736 6 right_width_0_height_0__pin_18_
port 24 nsew signal input
rlabel metal3 s 23800 11160 24600 11280 6 right_width_0_height_0__pin_19_
port 25 nsew signal input
rlabel metal3 s 23800 11704 24600 11824 6 right_width_0_height_0__pin_20_
port 26 nsew signal input
rlabel metal3 s 23800 12248 24600 12368 6 right_width_0_height_0__pin_21_
port 27 nsew signal input
rlabel metal3 s 23800 12792 24600 12912 6 right_width_0_height_0__pin_22_
port 28 nsew signal input
rlabel metal3 s 23800 13336 24600 13456 6 right_width_0_height_0__pin_23_
port 29 nsew signal input
rlabel metal3 s 23800 13880 24600 14000 6 right_width_0_height_0__pin_24_
port 30 nsew signal input
rlabel metal3 s 23800 14424 24600 14544 6 right_width_0_height_0__pin_25_
port 31 nsew signal input
rlabel metal3 s 23800 14968 24600 15088 6 right_width_0_height_0__pin_26_
port 32 nsew signal input
rlabel metal3 s 23800 15512 24600 15632 6 right_width_0_height_0__pin_27_
port 33 nsew signal input
rlabel metal3 s 23800 16056 24600 16176 6 right_width_0_height_0__pin_28_
port 34 nsew signal input
rlabel metal3 s 23800 16600 24600 16720 6 right_width_0_height_0__pin_29_
port 35 nsew signal input
rlabel metal3 s 23800 17144 24600 17264 6 right_width_0_height_0__pin_30_
port 36 nsew signal input
rlabel metal3 s 23800 17688 24600 17808 6 right_width_0_height_0__pin_31_
port 37 nsew signal input
rlabel metal3 s 23800 2456 24600 2576 6 right_width_0_height_0__pin_42_lower
port 38 nsew signal output
rlabel metal3 s 23800 18232 24600 18352 6 right_width_0_height_0__pin_42_upper
port 39 nsew signal output
rlabel metal3 s 23800 3000 24600 3120 6 right_width_0_height_0__pin_43_lower
port 40 nsew signal output
rlabel metal3 s 23800 18776 24600 18896 6 right_width_0_height_0__pin_43_upper
port 41 nsew signal output
rlabel metal3 s 23800 3544 24600 3664 6 right_width_0_height_0__pin_44_lower
port 42 nsew signal output
rlabel metal3 s 23800 19320 24600 19440 6 right_width_0_height_0__pin_44_upper
port 43 nsew signal output
rlabel metal3 s 23800 4088 24600 4208 6 right_width_0_height_0__pin_45_lower
port 44 nsew signal output
rlabel metal3 s 23800 19864 24600 19984 6 right_width_0_height_0__pin_45_upper
port 45 nsew signal output
rlabel metal3 s 23800 4632 24600 4752 6 right_width_0_height_0__pin_46_lower
port 46 nsew signal output
rlabel metal3 s 23800 20408 24600 20528 6 right_width_0_height_0__pin_46_upper
port 47 nsew signal output
rlabel metal3 s 23800 5176 24600 5296 6 right_width_0_height_0__pin_47_lower
port 48 nsew signal output
rlabel metal3 s 23800 20952 24600 21072 6 right_width_0_height_0__pin_47_upper
port 49 nsew signal output
rlabel metal3 s 23800 5720 24600 5840 6 right_width_0_height_0__pin_48_lower
port 50 nsew signal output
rlabel metal3 s 23800 21496 24600 21616 6 right_width_0_height_0__pin_48_upper
port 51 nsew signal output
rlabel metal3 s 23800 6264 24600 6384 6 right_width_0_height_0__pin_49_lower
port 52 nsew signal output
rlabel metal3 s 23800 22040 24600 22160 6 right_width_0_height_0__pin_49_upper
port 53 nsew signal output
rlabel metal2 s 5446 23800 5502 24600 6 top_width_0_height_0__pin_0_
port 54 nsew signal input
rlabel metal2 s 11886 23800 11942 24600 6 top_width_0_height_0__pin_10_
port 55 nsew signal input
rlabel metal2 s 12530 23800 12586 24600 6 top_width_0_height_0__pin_11_
port 56 nsew signal input
rlabel metal2 s 13174 23800 13230 24600 6 top_width_0_height_0__pin_12_
port 57 nsew signal input
rlabel metal2 s 13818 23800 13874 24600 6 top_width_0_height_0__pin_13_
port 58 nsew signal input
rlabel metal2 s 14462 23800 14518 24600 6 top_width_0_height_0__pin_14_
port 59 nsew signal input
rlabel metal2 s 15106 23800 15162 24600 6 top_width_0_height_0__pin_15_
port 60 nsew signal input
rlabel metal2 s 6090 23800 6146 24600 6 top_width_0_height_0__pin_1_
port 61 nsew signal input
rlabel metal2 s 6734 23800 6790 24600 6 top_width_0_height_0__pin_2_
port 62 nsew signal input
rlabel metal2 s 15750 23800 15806 24600 6 top_width_0_height_0__pin_32_
port 63 nsew signal input
rlabel metal2 s 16394 23800 16450 24600 6 top_width_0_height_0__pin_33_
port 64 nsew signal input
rlabel metal2 s 19614 23800 19670 24600 6 top_width_0_height_0__pin_34_lower
port 65 nsew signal output
rlabel metal2 s 294 23800 350 24600 6 top_width_0_height_0__pin_34_upper
port 66 nsew signal output
rlabel metal2 s 20258 23800 20314 24600 6 top_width_0_height_0__pin_35_lower
port 67 nsew signal output
rlabel metal2 s 938 23800 994 24600 6 top_width_0_height_0__pin_35_upper
port 68 nsew signal output
rlabel metal2 s 20902 23800 20958 24600 6 top_width_0_height_0__pin_36_lower
port 69 nsew signal output
rlabel metal2 s 1582 23800 1638 24600 6 top_width_0_height_0__pin_36_upper
port 70 nsew signal output
rlabel metal2 s 21546 23800 21602 24600 6 top_width_0_height_0__pin_37_lower
port 71 nsew signal output
rlabel metal2 s 2226 23800 2282 24600 6 top_width_0_height_0__pin_37_upper
port 72 nsew signal output
rlabel metal2 s 22190 23800 22246 24600 6 top_width_0_height_0__pin_38_lower
port 73 nsew signal output
rlabel metal2 s 2870 23800 2926 24600 6 top_width_0_height_0__pin_38_upper
port 74 nsew signal output
rlabel metal2 s 22834 23800 22890 24600 6 top_width_0_height_0__pin_39_lower
port 75 nsew signal output
rlabel metal2 s 3514 23800 3570 24600 6 top_width_0_height_0__pin_39_upper
port 76 nsew signal output
rlabel metal2 s 7378 23800 7434 24600 6 top_width_0_height_0__pin_3_
port 77 nsew signal input
rlabel metal2 s 23478 23800 23534 24600 6 top_width_0_height_0__pin_40_lower
port 78 nsew signal output
rlabel metal2 s 4158 23800 4214 24600 6 top_width_0_height_0__pin_40_upper
port 79 nsew signal output
rlabel metal2 s 24122 23800 24178 24600 6 top_width_0_height_0__pin_41_lower
port 80 nsew signal output
rlabel metal2 s 4802 23800 4858 24600 6 top_width_0_height_0__pin_41_upper
port 81 nsew signal output
rlabel metal2 s 8022 23800 8078 24600 6 top_width_0_height_0__pin_4_
port 82 nsew signal input
rlabel metal2 s 8666 23800 8722 24600 6 top_width_0_height_0__pin_5_
port 83 nsew signal input
rlabel metal2 s 9310 23800 9366 24600 6 top_width_0_height_0__pin_6_
port 84 nsew signal input
rlabel metal2 s 9954 23800 10010 24600 6 top_width_0_height_0__pin_7_
port 85 nsew signal input
rlabel metal2 s 10598 23800 10654 24600 6 top_width_0_height_0__pin_8_
port 86 nsew signal input
rlabel metal2 s 11242 23800 11298 24600 6 top_width_0_height_0__pin_9_
port 87 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 24600 24600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1873076
string GDS_FILE /home/marwan/clear_signoff_final/openlane/grid_clb/runs/grid_clb/results/signoff/grid_clb.magic.gds
string GDS_START 129632
<< end >>

