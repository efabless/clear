* NGSPICE file created from cby_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

.subckt cby_2__1_ IO_ISOL_N VGND VPWR ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ left_grid_pin_16_ left_grid_pin_17_ left_grid_pin_18_ left_grid_pin_19_ left_grid_pin_20_
+ left_grid_pin_21_ left_grid_pin_22_ left_grid_pin_23_ left_grid_pin_24_ left_grid_pin_25_
+ left_grid_pin_26_ left_grid_pin_27_ left_grid_pin_28_ left_grid_pin_29_ left_grid_pin_30_
+ left_grid_pin_31_ left_width_0_height_0__pin_0_ left_width_0_height_0__pin_1_lower
+ left_width_0_height_0__pin_1_upper prog_clk_0_N_out prog_clk_0_S_out prog_clk_0_W_in
+ right_grid_pin_0_
Xmux_right_ipin_11.mux_l2_in_0_ mux_right_ipin_11.mux_l1_in_1_/X mux_right_ipin_11.mux_l1_in_0_/X
+ mux_right_ipin_11.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_66_ _66_/A VGND VGND VPWR VPWR _66_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_11.mux_l1_in_1_ input35/X repeater119/X mux_right_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_49_ _49_/A VGND VGND VPWR VPWR _49_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput75 _72_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
Xoutput97 output97/A VGND VGND VPWR VPWR left_grid_pin_26_ sky130_fd_sc_hd__buf_2
Xoutput86 output86/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR sky130_fd_sc_hd__buf_2
Xoutput53 _50_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput64 _42_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_65_ _65_/A VGND VGND VPWR VPWR _65_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output95/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A0 _68_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_11.mux_l1_in_0_ input23/X repeater113/X mux_right_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_48_ _48_/A VGND VGND VPWR VPWR _48_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_0.mux_l2_in_3__130 VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/A0
+ mux_right_ipin_0.mux_l2_in_3__130/LO sky130_fd_sc_hd__conb_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput76 _73_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xoutput98 output98/A VGND VGND VPWR VPWR left_grid_pin_27_ sky130_fd_sc_hd__buf_2
XANTENNA_input30_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput87 output87/A VGND VGND VPWR VPWR left_grid_pin_16_ sky130_fd_sc_hd__buf_2
Xoutput54 _51_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput65 _43_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_7.mux_l2_in_3__126 VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/A0
+ mux_right_ipin_7.mux_l2_in_3__126/LO sky130_fd_sc_hd__conb_1
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_prog_clk_0_S_FTB01_A prog_clk_0_W_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_64_ _64_/A VGND VGND VPWR VPWR _64_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_3.mux_l2_in_3_ mux_right_ipin_3.mux_l2_in_3_/A0 _48_/A mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_3.mux_l2_in_2__A1 _42_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_47_ _47_/A VGND VGND VPWR VPWR _47_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_2.mux_l2_in_3__138 VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_3_/A0
+ mux_right_ipin_2.mux_l2_in_3__138/LO sky130_fd_sc_hd__conb_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_13.mux_l2_in_1__A0 _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_3.mux_l4_in_0_ mux_right_ipin_3.mux_l3_in_1_/X mux_right_ipin_3.mux_l3_in_0_/X
+ mux_right_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput66 _54_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput77 _55_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput99 output99/A VGND VGND VPWR VPWR left_grid_pin_28_ sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput55 _52_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xoutput88 output88/A VGND VGND VPWR VPWR left_grid_pin_17_ sky130_fd_sc_hd__buf_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_8.mux_l2_in_3_ mux_right_ipin_8.mux_l2_in_3_/A0 _53_/A mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l3_in_1_ mux_right_ipin_3.mux_l2_in_3_/X mux_right_ipin_3.mux_l2_in_2_/X
+ mux_right_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ _63_/A VGND VGND VPWR VPWR _63_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_3.mux_l2_in_2_ _68_/A _42_/A mux_right_ipin_3.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xprog_clk_0_FTB00 prog_clk_0_W_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmux_right_ipin_8.mux_l4_in_0_ mux_right_ipin_8.mux_l3_in_1_/X mux_right_ipin_8.mux_l3_in_0_/X
+ mux_right_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_46_ _46_/A VGND VGND VPWR VPWR _46_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_7.mux_l1_in_2__A0 _42_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l3_in_1_ mux_right_ipin_8.mux_l2_in_3_/X mux_right_ipin_8.mux_l2_in_2_/X
+ mux_right_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output88/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_11.mux_l2_in_3__A1 _50_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_1__A0 _66_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A0 _35_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput67 _64_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput78 _56_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_11.mux_l2_in_3__133 VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_3_/A0
+ mux_right_ipin_11.mux_l2_in_3__133/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput56 _53_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xoutput45 output45/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
Xoutput89 output89/A VGND VGND VPWR VPWR left_grid_pin_18_ sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_8.mux_l2_in_2_ _73_/A _47_/A mux_right_ipin_8.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input16_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.mux_l3_in_0_ mux_right_ipin_3.mux_l2_in_1_/X mux_right_ipin_3.mux_l2_in_0_/X
+ mux_right_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input8_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_62_ _62_/A VGND VGND VPWR VPWR _62_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_3.mux_l2_in_1_ _62_/A mux_right_ipin_3.mux_l1_in_2_/X mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_repeater118_A _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_45_ _45_/A VGND VGND VPWR VPWR _45_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_7.mux_l1_in_2__A1 _62_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l2_in_3_ mux_right_ipin_12.mux_l2_in_3_/A0 _51_/A mux_right_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l1_in_2_ _38_/A _58_/A mux_right_ipin_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_8.mux_l3_in_0_ mux_right_ipin_8.mux_l2_in_1_/X mux_right_ipin_8.mux_l2_in_0_/X
+ mux_right_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_10.mux_l1_in_0__A1 _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput46 _34_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput57 _35_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput68 _65_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xoutput79 _57_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_8.mux_l2_in_1_ _67_/A mux_right_ipin_8.mux_l1_in_2_/X mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_12.mux_l4_in_0_ mux_right_ipin_12.mux_l3_in_1_/X mux_right_ipin_12.mux_l3_in_0_/X
+ mux_right_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_5.mux_l2_in_3__A1 _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A0 _70_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l1_in_2_ _43_/A _63_/A mux_right_ipin_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_61_ _61_/A VGND VGND VPWR VPWR _61_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_12.mux_l3_in_1_ mux_right_ipin_12.mux_l2_in_3_/X mux_right_ipin_12.mux_l2_in_2_/X
+ mux_right_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_3.mux_l2_in_0_ mux_right_ipin_3.mux_l1_in_1_/X mux_right_ipin_3.mux_l1_in_0_/X
+ mux_right_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_44_ _44_/A VGND VGND VPWR VPWR _44_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input39_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l2_in_2_ _71_/A _47_/A mux_right_ipin_12.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_3.mux_l1_in_1_ _36_/A input15/X mux_right_ipin_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A0 _61_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput69 _66_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_8.mux_l2_in_0_ mux_right_ipin_8.mux_l1_in_1_/X mux_right_ipin_8.mux_l1_in_0_/X
+ mux_right_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput47 _44_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput58 _36_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input21_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_15.mux_l2_in_2__A1 _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_8.mux_l1_in_1_ repeater107/X repeater117/X mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_60_ _60_/A VGND VGND VPWR VPWR _60_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_12.mux_l3_in_0_ mux_right_ipin_12.mux_l2_in_1_/X mux_right_ipin_12.mux_l2_in_0_/X
+ mux_right_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__42__A _42_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__37__A _37_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A0 _68_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_43_ _43_/A VGND VGND VPWR VPWR _43_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_12.mux_l2_in_1_ _67_/A mux_right_ipin_12.mux_l1_in_2_/X mux_right_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_3.mux_l1_in_0_ _34_/A input3/X mux_right_ipin_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_2.mux_l2_in_1__A1 _37_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__50__A _50_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l1_in_2_ _41_/A _61_/A mux_right_ipin_12.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A0 _69_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput48 _45_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput59 _37_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__45__A _45_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_5.mux_l2_in_3__124 VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/A0
+ mux_right_ipin_5.mux_l2_in_3__124/LO sky130_fd_sc_hd__conb_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater120 input15/X VGND VGND VPWR VPWR _56_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input14_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_8.mux_l1_in_0_ repeater111/X repeater121/X mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input6_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR output86/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__53__A _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_9.mux_l2_in_2__A1 _40_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_42_ _42_/A VGND VGND VPWR VPWR _42_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output45_A output45/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l2_in_0_ mux_right_ipin_12.mux_l1_in_1_/X mux_right_ipin_12.mux_l1_in_0_/X
+ mux_right_ipin_12.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__48__A _48_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_12.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output99/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input44_A left_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_12.mux_l1_in_1_ repeater108/X repeater117/X mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output91/A sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_10.mux_l2_in_2__A1 _41_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput49 _46_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__61__A _61_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater110 input35/X VGND VGND VPWR VPWR repeater110/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater121 repeater122/X VGND VGND VPWR VPWR repeater121/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A0 _69_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_41_ _41_/A VGND VGND VPWR VPWR _41_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__64__A _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__59__A _59_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input37_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_12.mux_l1_in_0_ repeater112/X repeater121/X mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater111 repeater112/X VGND VGND VPWR VPWR repeater111/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater122 _55_/A VGND VGND VPWR VPWR repeater122/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__72__A _72_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_4.mux_l2_in_2__A1 _43_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_14.mux_l2_in_1__A0 _65_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_11.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_40_ _40_/A VGND VGND VPWR VPWR _40_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_4.mux_l2_in_3_ mux_right_ipin_4.mux_l2_in_3_/A0 _49_/A mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater112 _35_/A VGND VGND VPWR VPWR repeater112/X sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_ipin_0.mux_l2_in_3__129 VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_3_/A0
+ mux_left_ipin_0.mux_l2_in_3__129/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_4.mux_l4_in_0_ mux_right_ipin_4.mux_l3_in_1_/X mux_right_ipin_4.mux_l3_in_0_/X
+ mux_right_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_left_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_14.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_3_ mux_right_ipin_9.mux_l2_in_3_/A0 _48_/A mux_right_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l3_in_1_ mux_right_ipin_4.mux_l2_in_3_/X mux_right_ipin_4.mux_l2_in_2_/X
+ mux_right_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A0 _43_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_4.mux_l2_in_2_ _69_/A _43_/A mux_right_ipin_4.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.mux_l4_in_0_ mux_right_ipin_9.mux_l3_in_1_/X mux_right_ipin_9.mux_l3_in_0_/X
+ mux_right_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_3.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE input43/X
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR left_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_8
XANTENNA_input42_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l3_in_1_ mux_right_ipin_9.mux_l2_in_3_/X mux_right_ipin_9.mux_l2_in_2_/X
+ mux_right_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrepeater113 _54_/A VGND VGND VPWR VPWR repeater113/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_9.mux_l2_in_2_ _68_/A _40_/A mux_right_ipin_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l3_in_0_ mux_right_ipin_4.mux_l2_in_1_/X mux_right_ipin_4.mux_l2_in_0_/X
+ mux_right_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_8.mux_l1_in_2__A1 _63_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_4.mux_l2_in_1_ _63_/A mux_right_ipin_4.mux_l1_in_2_/X mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_15.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output102/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_13.mux_l2_in_3_ mux_right_ipin_13.mux_l2_in_3_/A0 _52_/A mux_right_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output94/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_4.mux_l1_in_2_ _39_/A _59_/A mux_right_ipin_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_6.mux_l2_in_3__A1 _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input35_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l3_in_0_ mux_right_ipin_9.mux_l2_in_1_/X mux_right_ipin_9.mux_l2_in_0_/X
+ mux_right_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater114 input3/X VGND VGND VPWR VPWR _54_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_3.mux_l1_in_2__A0 _38_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l2_in_1_ _60_/A repeater110/X mux_right_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_prog_clk_0_N_FTB01_A prog_clk_0_W_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_13.mux_l4_in_0_ mux_right_ipin_13.mux_l3_in_1_/X mux_right_ipin_13.mux_l3_in_0_/X
+ mux_right_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_3.mux_l2_in_1__A0 _62_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_13.mux_l3_in_1_ mux_right_ipin_13.mux_l2_in_3_/X mux_right_ipin_13.mux_l2_in_2_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l2_in_0_ mux_right_ipin_4.mux_l1_in_1_/X mux_right_ipin_4.mux_l1_in_0_/X
+ mux_right_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput1 IO_ISOL_N VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_13.mux_l2_in_2_ _72_/A _44_/A mux_right_ipin_13.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l1_in_1_ repeater107/X repeater118/X mux_right_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input28_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater115 repeater116/X VGND VGND VPWR VPWR _34_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xmem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_3.mux_l1_in_2__A1 _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_9.mux_l2_in_0_ _56_/A mux_right_ipin_9.mux_l1_in_0_/X mux_right_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_13.mux_l3_in_0_ mux_right_ipin_13.mux_l2_in_1_/X mux_right_ipin_13.mux_l2_in_0_/X
+ mux_right_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_3__A1 _48_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 ccff_head VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater112_A _35_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A0 _70_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_13.mux_l2_in_1_ _64_/A repeater110/X mux_right_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_4.mux_l1_in_0_ repeater111/X repeater122/X mux_right_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater116 input23/X VGND VGND VPWR VPWR repeater116/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_ipin_0.mux_l2_in_3__A1 _50_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input40_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output87/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_14.mux_l2_in_3__136 VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/A0
+ mux_right_ipin_14.mux_l2_in_3__136/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_9.mux_l1_in_0_ repeater116/X _54_/A mux_right_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chany_bottom_in[0] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_11.mux_l2_in_2__A1 _46_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_13.mux_l2_in_0_ repeater119/X mux_right_ipin_13.mux_l1_in_0_/X mux_right_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater117 repeater118/X VGND VGND VPWR VPWR repeater117/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_W_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input33_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A0 _72_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 chany_bottom_in[10] VGND VGND VPWR VPWR _64_/A sky130_fd_sc_hd__clkbuf_2
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_15.mux_l1_in_2__A0 _38_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput40 chany_top_in[7] VGND VGND VPWR VPWR _41_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater107 repeater108/X VGND VGND VPWR VPWR repeater107/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater118 _57_/A VGND VGND VPWR VPWR repeater118/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input26_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_2__A1 _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_13.mux_l1_in_0_ repeater116/X repeater113/X mux_right_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_15.mux_l2_in_1__A0 _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l2_in_3_ mux_right_ipin_0.mux_l2_in_3_/A0 _51_/A mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_2.mux_l2_in_0__A0 _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 chany_bottom_in[11] VGND VGND VPWR VPWR _65_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ mux_right_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_59_ _59_/A VGND VGND VPWR VPWR _59_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_15.mux_l1_in_2__A1 _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_5.mux_l2_in_3_ mux_right_ipin_5.mux_l2_in_3_/A0 _52_/A mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l2_in_3__131 VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_3_/A0
+ mux_right_ipin_1.mux_l2_in_3__131/LO sky130_fd_sc_hd__conb_1
Xinput41 chany_top_in[8] VGND VGND VPWR VPWR _42_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater108 _37_/A VGND VGND VPWR VPWR repeater108/X sky130_fd_sc_hd__clkbuf_1
Xrepeater119 _56_/A VGND VGND VPWR VPWR repeater119/X sky130_fd_sc_hd__clkbuf_1
Xinput30 chany_top_in[16] VGND VGND VPWR VPWR _50_/A sky130_fd_sc_hd__clkbuf_2
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input19_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_0.mux_l2_in_2_ _71_/A _45_/A mux_right_ipin_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l4_in_0_ mux_right_ipin_5.mux_l3_in_1_/X mux_right_ipin_5.mux_l3_in_0_/X
+ mux_right_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_13.mux_l2_in_3__A1 _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_8.mux_l2_in_3__127 VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/A0
+ mux_right_ipin_8.mux_l2_in_3__127/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_9.mux_l2_in_1__A0 _60_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l3_in_1_ mux_right_ipin_5.mux_l2_in_3_/X mux_right_ipin_5.mux_l2_in_2_/X
+ mux_right_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 chany_bottom_in[12] VGND VGND VPWR VPWR _66_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__40__A _40_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_58_ _58_/A VGND VGND VPWR VPWR _58_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_0.mux_l2_in_2__A1 _45_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A0 _61_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_5.mux_l2_in_2_ _72_/A _44_/A mux_right_ipin_5.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__35__A _35_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.mux_l2_in_3__139 VGND VGND VPWR VPWR mux_right_ipin_3.mux_l2_in_3_/A0
+ mux_right_ipin_3.mux_l2_in_3__139/LO sky130_fd_sc_hd__conb_1
Xinput31 chany_top_in[17] VGND VGND VPWR VPWR _51_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrepeater109 repeater110/X VGND VGND VPWR VPWR _36_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chany_bottom_in[7] VGND VGND VPWR VPWR _61_/A sky130_fd_sc_hd__clkbuf_2
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput42 chany_top_in[9] VGND VGND VPWR VPWR _43_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_11.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output98/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input31_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l2_in_1_ _65_/A mux_right_ipin_0.mux_l1_in_2_/X mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output90/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__43__A _43_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l1_in_2_ _39_/A _59_/A mux_right_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_5.mux_l3_in_0_ mux_right_ipin_5.mux_l2_in_1_/X mux_right_ipin_5.mux_l2_in_0_/X
+ mux_right_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__38__A _38_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_74_ left_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR _74_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_7.mux_l2_in_3__A1 _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chany_bottom_in[13] VGND VGND VPWR VPWR _67_/A sky130_fd_sc_hd__clkbuf_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_57_ _57_/A VGND VGND VPWR VPWR _57_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_5.mux_l2_in_1_ _64_/A _36_/A mux_right_ipin_5.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_10.mux_l2_in_1__A1 _37_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A0 _39_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput32 chany_top_in[18] VGND VGND VPWR VPWR _52_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 gfpga_pad_EMBEDDED_IO_HD_SOC_IN VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput10 chany_bottom_in[16] VGND VGND VPWR VPWR _70_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 chany_bottom_in[8] VGND VGND VPWR VPWR _62_/A sky130_fd_sc_hd__clkbuf_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE input44/X
+ output86/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT sky130_fd_sc_hd__ebufn_8
XANTENNA__46__A _46_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l2_in_3_ mux_right_ipin_14.mux_l2_in_3_/A0 _53_/A mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l2_in_1__A0 _63_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input24_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_12.mux_l2_in_3__134 VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_3_/A0
+ mux_right_ipin_12.mux_l2_in_3__134/LO sky130_fd_sc_hd__conb_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.mux_l4_in_0_ mux_right_ipin_14.mux_l3_in_1_/X mux_right_ipin_14.mux_l3_in_0_/X
+ mux_right_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_0.mux_l1_in_1_ repeater107/X repeater118/X mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_73_ _73_/A VGND VGND VPWR VPWR _73_/X sky130_fd_sc_hd__clkbuf_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 chany_bottom_in[14] VGND VGND VPWR VPWR _68_/A sky130_fd_sc_hd__clkbuf_2
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__49__A _49_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_56_ _56_/A VGND VGND VPWR VPWR _56_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_14.mux_l3_in_1_ mux_right_ipin_14.mux_l2_in_3_/X mux_right_ipin_14.mux_l2_in_2_/X
+ mux_right_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_5.mux_l2_in_0_ input15/X mux_right_ipin_5.mux_l1_in_0_/X mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_4.mux_l1_in_2__A1 _59_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput33 chany_top_in[19] VGND VGND VPWR VPWR _53_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 left_width_0_height_0__pin_0_ VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
X_39_ _39_/A VGND VGND VPWR VPWR _39_/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chany_bottom_in[9] VGND VGND VPWR VPWR _63_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chany_bottom_in[17] VGND VGND VPWR VPWR _71_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__62__A _62_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l2_in_2_ _73_/A _45_/A mux_right_ipin_14.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__57__A _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input17_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_2.mux_l2_in_3__A1 _49_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_0.mux_l1_in_0_ repeater111/X repeater122/X mux_right_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__70__A _70_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ _72_/A VGND VGND VPWR VPWR _72_/X sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 chany_bottom_in[15] VGND VGND VPWR VPWR _69_/A sky130_fd_sc_hd__clkbuf_2
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__65__A _65_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_55_ _55_/A VGND VGND VPWR VPWR _55_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_14.mux_l3_in_0_ mux_right_ipin_14.mux_l2_in_1_/X mux_right_ipin_14.mux_l2_in_0_/X
+ mux_right_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput34 chany_top_in[1] VGND VGND VPWR VPWR _35_/A sky130_fd_sc_hd__clkbuf_2
Xinput23 chany_top_in[0] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput12 chany_bottom_in[18] VGND VGND VPWR VPWR _72_/A sky130_fd_sc_hd__clkbuf_2
X_38_ _38_/A VGND VGND VPWR VPWR _38_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_ipin_14.mux_l2_in_1_ _65_/A repeater108/X mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_5.mux_l1_in_0_ _34_/A input3/X mux_right_ipin_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A _68_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_71_ _71_/A VGND VGND VPWR VPWR _71_/X sky130_fd_sc_hd__clkbuf_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_54_ _54_/A VGND VGND VPWR VPWR _54_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xoutput100 output100/A VGND VGND VPWR VPWR left_grid_pin_29_ sky130_fd_sc_hd__buf_2
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xinput24 chany_top_in[10] VGND VGND VPWR VPWR _44_/A sky130_fd_sc_hd__clkbuf_2
Xinput35 chany_top_in[2] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 chany_bottom_in[19] VGND VGND VPWR VPWR _73_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_37_ _37_/A VGND VGND VPWR VPWR _37_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_14.mux_l2_in_0_ repeater117/X mux_right_ipin_14.mux_l1_in_0_/X mux_right_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_14.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output101/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_6.mux_l2_in_3__125 VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_3_/A0
+ mux_right_ipin_6.mux_l2_in_3__125/LO sky130_fd_sc_hd__conb_1
XANTENNA_input22_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output93/A sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_70_ _70_/A VGND VGND VPWR VPWR _70_/X sky130_fd_sc_hd__clkbuf_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_53_ _53_/A VGND VGND VPWR VPWR _53_/X sky130_fd_sc_hd__clkbuf_1
Xoutput101 output101/A VGND VGND VPWR VPWR left_grid_pin_30_ sky130_fd_sc_hd__buf_2
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_6.mux_l2_in_2__A1 _45_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput36 chany_top_in[3] VGND VGND VPWR VPWR _37_/A sky130_fd_sc_hd__clkbuf_2
Xinput25 chany_top_in[11] VGND VGND VPWR VPWR _45_/A sky130_fd_sc_hd__clkbuf_2
Xinput14 chany_bottom_in[1] VGND VGND VPWR VPWR _55_/A sky130_fd_sc_hd__clkbuf_2
X_36_ _36_/A VGND VGND VPWR VPWR _36_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_5.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_14.mux_l1_in_0_ repeater112/X repeater121/X mux_right_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input15_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input7_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.mux_l2_in_3_ mux_right_ipin_1.mux_l2_in_3_/A0 _48_/A mux_right_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A0 _68_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ _52_/A VGND VGND VPWR VPWR _52_/X sky130_fd_sc_hd__clkbuf_1
Xoutput102 output102/A VGND VGND VPWR VPWR left_grid_pin_31_ sky130_fd_sc_hd__buf_2
Xmem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput26 chany_top_in[12] VGND VGND VPWR VPWR _46_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 chany_top_in[4] VGND VGND VPWR VPWR _38_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xmux_right_ipin_1.mux_l4_in_0_ mux_right_ipin_1.mux_l3_in_1_/X mux_right_ipin_1.mux_l3_in_0_/X
+ mux_right_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_35_ _35_/A VGND VGND VPWR VPWR _35_/X sky130_fd_sc_hd__clkbuf_1
Xinput15 chany_bottom_in[2] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A0 _70_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X mux_right_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR output45/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_14.mux_l2_in_3__A1 _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_6.mux_l2_in_3_ mux_right_ipin_6.mux_l2_in_3_/A0 _53_/A mux_right_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l3_in_1_ mux_right_ipin_1.mux_l2_in_3_/X mux_right_ipin_1.mux_l2_in_2_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_10.mux_l2_in_3__132 VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/A0
+ mux_right_ipin_10.mux_l2_in_3__132/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_11.mux_l1_in_2__A0 _40_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_left_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_1.mux_l2_in_2_ _68_/A _40_/A mux_right_ipin_1.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_ipin_1.mux_l2_in_2__A1 _40_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_6.mux_l4_in_0_ mux_right_ipin_6.mux_l3_in_1_/X mux_right_ipin_6.mux_l3_in_0_/X
+ mux_right_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_11.mux_l2_in_1__A0 _66_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_13.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput103 _74_/X VGND VGND VPWR VPWR left_width_0_height_0__pin_1_upper sky130_fd_sc_hd__buf_2
X_51_ _51_/A VGND VGND VPWR VPWR _51_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_0_S_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR output105/A sky130_fd_sc_hd__buf_4
Xmux_right_ipin_6.mux_l3_in_1_ mux_right_ipin_6.mux_l2_in_3_/X mux_right_ipin_6.mux_l2_in_2_/X
+ mux_right_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput27 chany_top_in[13] VGND VGND VPWR VPWR _47_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 chany_top_in[5] VGND VGND VPWR VPWR _39_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 chany_bottom_in[3] VGND VGND VPWR VPWR _57_/A sky130_fd_sc_hd__clkbuf_2
X_34_ _34_/A VGND VGND VPWR VPWR _34_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_ipin_0.mux_l2_in_2__A1 _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input38_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_6.mux_l2_in_2_ _73_/A _45_/A mux_right_ipin_6.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_1.mux_l3_in_0_ mux_right_ipin_1.mux_l2_in_1_/X mux_right_ipin_1.mux_l2_in_0_/X
+ mux_right_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_11.mux_l1_in_2__A1 _60_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_8.mux_l2_in_3__A1 _53_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_1.mux_l2_in_1_ _60_/A repeater110/X mux_right_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput104 output104/A VGND VGND VPWR VPWR prog_clk_0_N_out sky130_fd_sc_hd__clkbuf_1
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_A
+ output45/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_50_ _50_/A VGND VGND VPWR VPWR _50_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_10.mux_l2_in_3_ mux_right_ipin_10.mux_l2_in_3_/A0 _49_/A mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l3_in_0_ mux_right_ipin_6.mux_l2_in_1_/X mux_right_ipin_6.mux_l2_in_0_/X
+ mux_right_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput39 chany_top_in[6] VGND VGND VPWR VPWR _40_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 chany_top_in[14] VGND VGND VPWR VPWR _48_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput17 chany_bottom_in[4] VGND VGND VPWR VPWR _58_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater122_A _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_5.mux_l2_in_1__A0 _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_6.mux_l2_in_1_ _65_/A repeater107/X mux_right_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_10.mux_l4_in_0_ mux_right_ipin_10.mux_l3_in_1_/X mux_right_ipin_10.mux_l3_in_0_/X
+ mux_right_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l2_in_3_ mux_right_ipin_15.mux_l2_in_3_/A0 _50_/A mux_right_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_left_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_10.mux_l3_in_1_ mux_right_ipin_10.mux_l2_in_3_/X mux_right_ipin_10.mux_l2_in_2_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output96/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_1.mux_l2_in_0_ _56_/A mux_right_ipin_1.mux_l1_in_0_/X mux_right_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input13_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_10.mux_l2_in_2_ _69_/A _41_/A mux_right_ipin_10.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput105 output105/A VGND VGND VPWR VPWR prog_clk_0_S_out sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_15.mux_l4_in_0_ mux_right_ipin_15.mux_l3_in_1_/X mux_right_ipin_15.mux_l3_in_0_/X
+ mux_right_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput29 chany_top_in[15] VGND VGND VPWR VPWR _49_/A sky130_fd_sc_hd__clkbuf_2
Xinput18 chany_bottom_in[5] VGND VGND VPWR VPWR _59_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_ipin_15.mux_l3_in_1_ mux_right_ipin_15.mux_l2_in_3_/X mux_right_ipin_15.mux_l2_in_2_/X
+ mux_right_ipin_15.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_6.mux_l2_in_0_ repeater117/X mux_right_ipin_6.mux_l1_in_0_/X mux_right_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input43_A gfpga_pad_EMBEDDED_IO_HD_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_3.mux_l2_in_3__A1 _48_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A0 _35_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_4.mux_l2_in_3__123 VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/A0
+ mux_right_ipin_4.mux_l2_in_3__123/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A0 _72_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l2_in_2_ _70_/A _44_/A mux_right_ipin_15.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X input2/X VGND VGND
+ VPWR VPWR mux_left_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_10.mux_l3_in_0_ mux_right_ipin_10.mux_l2_in_1_/X mux_right_ipin_10.mux_l2_in_0_/X
+ mux_right_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A0 _39_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_0.mux_l2_in_1__A0 _65_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_10.mux_l2_in_1_ _61_/A _37_/A mux_right_ipin_10.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_1.mux_l1_in_0_ repeater116/X _54_/A mux_right_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput106 output106/A VGND VGND VPWR VPWR right_grid_pin_0_ sky130_fd_sc_hd__buf_2
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 chany_bottom_in[6] VGND VGND VPWR VPWR _60_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater108_A _37_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_15.mux_l3_in_0_ mux_right_ipin_15.mux_l2_in_1_/X mux_right_ipin_15.mux_l2_in_0_/X
+ mux_right_ipin_15.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_ipin_2.mux_l1_in_0__A1 _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_13.mux_l2_in_2__A1 _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l2_in_1_ _64_/A mux_right_ipin_15.mux_l1_in_2_/X mux_right_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l2_in_3_ mux_left_ipin_0.mux_l2_in_3_/A0 _50_/A mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_6.mux_l1_in_0_ repeater111/X repeater121/X mux_right_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_0.mux_l1_in_2__A1 _59_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A0 _72_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_15.mux_l1_in_2_ _38_/A _58_/A mux_right_ipin_15.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l2_in_0_ _57_/A mux_right_ipin_10.mux_l1_in_0_/X mux_right_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_10.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output97/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_ipin_10.mux_l2_in_0__A0 _57_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l4_in_0_ mux_left_ipin_0.mux_l3_in_1_/X mux_left_ipin_0.mux_l3_in_0_/X
+ mux_left_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output89/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_ipin_0.mux_l3_in_1_ mux_left_ipin_0.mux_l2_in_3_/X mux_left_ipin_0.mux_l2_in_2_/X
+ mux_left_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input29_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_15.mux_l2_in_0_ mux_right_ipin_15.mux_l1_in_1_/X mux_right_ipin_15.mux_l1_in_0_/X
+ mux_right_ipin_15.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l2_in_2_ _70_/A _44_/A mux_left_ipin_0.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR mux_left_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_1_ input35/X repeater119/X mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_7.mux_l2_in_2__A1 _46_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l2_in_3__137 VGND VGND VPWR VPWR mux_right_ipin_15.mux_l2_in_3_/A0
+ mux_right_ipin_15.mux_l2_in_3__137/LO sky130_fd_sc_hd__conb_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput90 output90/A VGND VGND VPWR VPWR left_grid_pin_19_ sky130_fd_sc_hd__buf_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input3_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__41__A _41_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_10.mux_l1_in_0_ _35_/A _55_/A mux_right_ipin_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_right_ipin_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_ipin_0.mux_l3_in_0_ mux_left_ipin_0.mux_l2_in_1_/X mux_left_ipin_0.mux_l2_in_0_/X
+ mux_left_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input41_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A0 _69_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.mux_l2_in_1_ _64_/A mux_left_ipin_0.mux_l1_in_2_/X mux_left_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__44__A _44_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_ipin_15.mux_l1_in_0_ input23/X repeater113/X mux_right_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_ipin_0.mux_l1_in_2_ _38_/A _58_/A mux_left_ipin_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR mux_left_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__39__A _39_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput80 _58_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_2.mux_l2_in_3_ mux_right_ipin_2.mux_l2_in_3_/A0 _49_/A mux_right_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xoutput91 output91/A VGND VGND VPWR VPWR left_grid_pin_20_ sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_ipin_15.mux_l2_in_3__A1 _50_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__52__A _52_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_N_FTB01 prog_clk_0_W_in VGND VGND VPWR VPWR output104/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A0 _41_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l4_in_0_ mux_right_ipin_2.mux_l3_in_1_/X mux_right_ipin_2.mux_l3_in_0_/X
+ mux_right_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_2__A1 _41_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input34_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_7.mux_l2_in_3_ mux_right_ipin_7.mux_l2_in_3_/A0 _52_/A mux_right_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_ipin_0.mux_l2_in_0_ mux_left_ipin_0.mux_l1_in_1_/X mux_left_ipin_0.mux_l1_in_0_/X
+ mux_left_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_2.mux_l3_in_1_ mux_right_ipin_2.mux_l2_in_3_/X mux_right_ipin_2.mux_l2_in_2_/X
+ mux_right_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__60__A _60_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__55__A _55_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_ipin_0.mux_l1_in_1_ _36_/A input15/X mux_left_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput70 _67_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput81 _59_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput92 output92/A VGND VGND VPWR VPWR left_grid_pin_21_ sky130_fd_sc_hd__buf_2
Xmux_right_ipin_7.mux_l4_in_0_ mux_right_ipin_7.mux_l3_in_1_/X mux_right_ipin_7.mux_l3_in_0_/X
+ mux_right_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_ipin_2.mux_l2_in_2_ _69_/A _41_/A mux_right_ipin_2.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE output45/A
+ input1/X VGND VGND VPWR VPWR output86/A sky130_fd_sc_hd__or2b_2
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_7.mux_l3_in_1_ mux_right_ipin_7.mux_l2_in_3_/X mux_right_ipin_7.mux_l2_in_2_/X
+ mux_right_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__63__A _63_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_ipin_12.mux_l1_in_2__A1 _61_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_9.mux_l2_in_3__A1 _48_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__58__A _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_7.mux_l2_in_2_ _72_/A _46_/A mux_right_ipin_7.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_7.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_2.mux_l3_in_0_ mux_right_ipin_2.mux_l2_in_1_/X mux_right_ipin_2.mux_l2_in_0_/X
+ mux_right_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_ipin_10.mux_l2_in_3__A1 _49_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_ipin_0.mux_l1_in_0_ _34_/A input3/X mux_left_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput71 _68_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xoutput82 _60_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_9.mux_l2_in_3__128 VGND VGND VPWR VPWR mux_right_ipin_9.mux_l2_in_3_/A0
+ mux_right_ipin_9.mux_l2_in_3__128/LO sky130_fd_sc_hd__conb_1
Xoutput93 output93/A VGND VGND VPWR VPWR left_grid_pin_22_ sky130_fd_sc_hd__buf_2
Xoutput60 _38_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_2.mux_l2_in_1_ _61_/A _37_/A mux_right_ipin_2.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_ipin_6.mux_l2_in_1__A0 _65_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_13.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR output100/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__66__A _66_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output92/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input1_A IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_11.mux_l2_in_3_ mux_right_ipin_11.mux_l2_in_3_/A0 _50_/A mux_right_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_69_ _69_/A VGND VGND VPWR VPWR _69_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_7.mux_l3_in_0_ mux_right_ipin_7.mux_l2_in_1_/X mux_right_ipin_7.mux_l2_in_0_/X
+ mux_right_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__74__A left_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_12.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l2_in_1_ _66_/A mux_right_ipin_7.mux_l1_in_2_/X mux_right_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__69__A _69_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l4_in_0_ mux_right_ipin_11.mux_l3_in_1_/X mux_right_ipin_11.mux_l3_in_0_/X
+ mux_right_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput72 _69_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput83 _61_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_7.mux_l1_in_2_ _42_/A _62_/A mux_right_ipin_7.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput94 output94/A VGND VGND VPWR VPWR left_grid_pin_23_ sky130_fd_sc_hd__buf_2
Xoutput50 _47_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput61 _39_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_11.mux_l3_in_1_ mux_right_ipin_11.mux_l2_in_3_/X mux_right_ipin_11.mux_l2_in_2_/X
+ mux_right_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_2.mux_l2_in_0_ _57_/A mux_right_ipin_2.mux_l1_in_0_/X mux_right_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_2.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_left_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output106/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_ipin_4.mux_l2_in_3__A1 _49_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l2_in_2_ _70_/A _46_/A mux_right_ipin_11.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_68_ _68_/A VGND VGND VPWR VPWR _68_/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_right_ipin_15.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_1.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l2_in_0_ mux_right_ipin_7.mux_l1_in_1_/X mux_right_ipin_7.mux_l1_in_0_/X
+ mux_right_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input32_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_ipin_1.mux_l2_in_1__A0 _60_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput73 _70_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xoutput84 _62_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xmux_right_ipin_13.mux_l2_in_3__135 VGND VGND VPWR VPWR mux_right_ipin_13.mux_l2_in_3_/A0
+ mux_right_ipin_13.mux_l2_in_3__135/LO sky130_fd_sc_hd__conb_1
Xmux_right_ipin_7.mux_l1_in_1_ input35/X repeater119/X mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput95 output95/A VGND VGND VPWR VPWR left_grid_pin_24_ sky130_fd_sc_hd__buf_2
Xoutput51 _48_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput62 _40_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A0 _38_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l3_in_0_ mux_right_ipin_11.mux_l2_in_1_/X mux_right_ipin_11.mux_l2_in_0_/X
+ mux_right_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_4.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_ipin_0.mux_l2_in_1__A0 _64_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_11.mux_l2_in_1_ _66_/A mux_right_ipin_11.mux_l1_in_2_/X mux_right_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_2.mux_l1_in_0_ _35_/A _55_/A mux_right_ipin_2.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_right_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_67_ _67_/A VGND VGND VPWR VPWR _67_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_ipin_14.mux_l2_in_2__A1 _45_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_right_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_15.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_11.mux_l1_in_2_ _40_/A _60_/A mux_right_ipin_11.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_11.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_right_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_12.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input25_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_right_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_ipin_7.mux_l1_in_0_ input23/X repeater113/X mux_right_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput52 _49_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_ipin_0.mux_l1_in_2__A1 _58_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput74 _71_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput85 _63_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput96 output96/A VGND VGND VPWR VPWR left_grid_pin_25_ sky130_fd_sc_hd__buf_2
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 _41_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
.ends

