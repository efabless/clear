* NGSPICE file created from bottom_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

.subckt bottom_tile VGND VPWR ccff_head ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0]
+ chanx_right_in_0[10] chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13]
+ chanx_right_in_0[14] chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17]
+ chanx_right_in_0[18] chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20]
+ chanx_right_in_0[21] chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24]
+ chanx_right_in_0[25] chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28]
+ chanx_right_in_0[29] chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4]
+ chanx_right_in_0[5] chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8]
+ chanx_right_in_0[9] chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11]
+ chanx_right_out_0[12] chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15]
+ chanx_right_out_0[16] chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19]
+ chanx_right_out_0[1] chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22]
+ chanx_right_out_0[23] chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26]
+ chanx_right_out_0[27] chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2]
+ chanx_right_out_0[3] chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6]
+ chanx_right_out_0[7] chanx_right_out_0[8] chanx_right_out_0[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[20] chany_top_in[21] chany_top_in[22] chany_top_in[23] chany_top_in[24]
+ chany_top_in[25] chany_top_in[26] chany_top_in[27] chany_top_in[28] chany_top_in[29]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[20] chany_top_out[21] chany_top_out[22] chany_top_out[23] chany_top_out[24]
+ chany_top_out[25] chany_top_out[26] chany_top_out[27] chany_top_out[28] chany_top_out[29]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1]
+ gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1]
+ gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1]
+ gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset reset
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
+ top_width_0_height_0_subtile_0__pin_inpad_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ top_width_0_height_0_subtile_2__pin_inpad_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold340 sb_1__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold351 sb_1__0_.mem_top_track_4.mem_out\[0\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold362 sb_1__0_.mem_right_track_52.mem_out\[0\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold384 net417 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold373 sb_1__0_.mem_right_track_10.mem_out\[0\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_hold374_A sb_1__0_.mem_top_track_8.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net344
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_input92_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_29.mux_l1_in_1_ net39 net86 sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_40.mux_l2_in_0__250 VGND VGND VPWR VPWR net250 sb_1__0_.mux_top_track_40.mux_l2_in_0__250/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 net278 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold181 sb_1__0_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold192 net289 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mux_right_track_0.mux_l1_in_0_ net91 net73 sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net519
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_4.mux_l2_in_1_ net249 net17 sb_1__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net541
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__124__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_ net260 net58 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__S sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__S sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk net437
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net467
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
X_131_ sb_1__0_.mux_left_track_5.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk net493
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input55_A chanx_right_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__119__A sb_1__0_.mux_left_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_28.mux_l1_in_0_ net29 net59 sb_1__0_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_30.mux_l1_in_0_ net28 net58 sb_1__0_.mem_top_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l3_in_0__S sb_1__0_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_ net35 net4 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__S sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_114_ net35 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_42.mux_l2_in_0_ net251 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0 net39 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net407
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xhold74 net538 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 net464 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 net478 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold63 net526 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold41 net542 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold96 net599 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold85 net570 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_5 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout205_A net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__127__A sb_1__0_.mux_left_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_58.mux_l2_in_0__S sb_1__0_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__S sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xhold363 sb_1__0_.mem_top_track_0.mem_out\[1\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold374 sb_1__0_.mem_top_track_8.mem_out\[0\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold330 sb_1__0_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold385 net2 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold352 sb_1__0_.mem_top_track_16.mem_out\[1\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold341 sb_1__0_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net547
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input85_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l1_in_0_ net68 net80 sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold182 net284 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold171 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold193 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold160 net273 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net497
+ net215 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_4.mux_l2_in_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__140__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_ net27 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_22.mux_l1_in_1__241 VGND VGND VPWR VPWR net241 sb_1__0_.mux_top_track_22.mux_l1_in_1__241/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_130_ sb_1__0_.mux_left_track_7.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chanx_right_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__135__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_4.mux_l1_in_1_ net47 net50 sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input102_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ net34 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_ net41 net10 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net463
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold86 net568 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold64 net528 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold97 net596 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 net456 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 net556 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold31 net482 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 net486 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 net484 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 net252 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_18.mux_l2_in_1__238 VGND VGND VPWR VPWR net238 sb_1__0_.mux_top_track_18.mux_l2_in_1__238/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_42.mux_l1_in_0_ net27 net100 sb_1__0_.mem_top_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__143__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.out sky130_fd_sc_hd__clkbuf_1
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold320 sb_1__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold342 sb_1__0_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold364 sb_1__0_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold331 sb_1__0_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold375 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net642
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold386 ccff_head VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold353 sb_1__0_.mem_right_track_36.mem_out\[0\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input78_A chany_top_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__138__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold183 sb_1__0_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold150 net650 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold172 net280 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold161 sb_1__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold194 net292 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput200 net200 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_189_ sb_1__0_.mux_top_track_8.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__151__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_4.mux_l1_in_0_ net102 net99 sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_28.mux_l3_in_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold342_A sb_1__0_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_112_ net62 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__146__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l2_in_0__S sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_45.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A1 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xhold98 net593 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold10 net434 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_2
Xhold76 net581 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold43 net532 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 net476 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 net450 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 net488 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold65 net546 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold87 net585 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ net372 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l2_in_1_ net227 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_28.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput100 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net527
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__S sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold310 net351 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_fanout210_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold321 net356 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold332 sb_1__0_.mem_top_track_10.mem_out\[0\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold343 sb_1__0_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold354 sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold376 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net643
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold365 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net632
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold387 net420 VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_28.mux_l1_in_2_ net14 net9 sb_1__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__154__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net375
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold140 net637 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold151 net652 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold162 net275 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold195 sb_1__0_.mem_right_track_0.ccff_tail VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold184 net288 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold173 sb_1__0_.mem_top_track_36.ccff_tail VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold372_A sb_1__0_.mem_top_track_2.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_12.mux_l3_in_0_ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input90_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput201 net201 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_9_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_0.mux_l1_in_3__233 VGND VGND VPWR VPWR net233 sb_1__0_.mux_top_track_0.mux_l1_in_3__233/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__S sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_188_ sb_1__0_.mux_top_track_10.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_53.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ net579 net207 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_top_track_12.mux_l2_in_1_ net235 net11 sb_1__0_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_18_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold168_A net277 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_20.mux_l2_in_1__226 VGND VGND VPWR VPWR net226 sb_1__0_.mux_right_track_20.mux_l2_in_1__226/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_111_ sb_1__0_.mux_left_track_45.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_2_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_45.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 net436 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold22 net458 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold55 net540 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 net480 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold66 net558 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold88 net589 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold77 net586 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold99 net600 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 net518 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ net358 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_28.mux_l2_in_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net101 sky130_fd_sc_hd__buf_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net571
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_13.mux_l3_in_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold322 sb_1__0_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_fanout203_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold311 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net578
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold344 sb_1__0_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold300 net346 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold333 sb_1__0_.mem_right_track_10.mem_out\[1\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold355 sb_1__0_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold377 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net644
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold366 sb_1__0_.mem_top_track_18.mem_out\[1\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold388 net270 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ net74 sb_1__0_.mem_right_track_28.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net394
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold163 sb_1__0_.mem_top_track_10.ccff_tail VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold152 net269 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold185 sb_1__0_.mem_top_track_42.mem_out\[0\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold141 net642 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold174 net276 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold130 net623 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_left_track_13.mux_l2_in_1_ net265 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xhold196 net291 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input83_A chany_top_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput202 net202 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_9_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_187_ sb_1__0_.mux_top_track_12.out VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_left_track_53.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ net405 net207 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_12.mux_l2_in_0_ net36 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_13.mux_l1_in_2_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net56 sb_1__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_52.mux_l1_in_1__231 VGND VGND VPWR VPWR net231 sb_1__0_.mux_right_track_52.mux_l1_in_1__231/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ net60 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_ sb_1__0_.mux_left_track_3.out net23
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input46_A chanx_right_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold45 net504 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold34 net472 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 net500 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold12 net444 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 net468 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold78 net574 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold89 net587 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input100_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold67 net544 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_9 net253 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net412 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
+ clknet_4_2_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_11.mux_l1_in_3__264 VGND VGND VPWR VPWR net264 sb_1__0_.mux_left_track_11.mux_l1_in_3__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net102 sky130_fd_sc_hd__buf_2
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_50.mux_l2_in_0__A0 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__S sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold345 sb_1__0_.mem_top_track_6.mem_out\[0\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold301 sb_1__0_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold334 sb_1__0_.mem_top_track_8.mem_out\[1\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold323 sb_1__0_.mem_right_track_20.mem_out\[0\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold378 sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold312 net347 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold356 sb_1__0_.mem_top_track_36.mem_out\[0\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0 sb_1__0_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold367 sb_1__0_.mem_right_track_28.mem_out\[0\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold389 net421 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l1_in_0_ net66 net78 sb_1__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net354
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk net327
+ net208 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_6.mux_l1_in_3_ net232 net29 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold142 net639 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold164 net281 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold186 net286 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold197 sb_1__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold120 net614 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold153 net653 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold131 net628 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__261 VGND VGND VPWR VPWR net261 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__261/LO
+ sky130_fd_sc_hd__conb_1
Xhold175 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__S sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_13.mux_l2_in_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold358_A sb_1__0_.mem_right_track_6.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input76_A chany_top_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_50.mux_l2_in_0__S sb_1__0_.mem_top_track_50.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__S sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_186_ sb_1__0_.mux_top_track_14.out VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_0_0_prog_clk net423 net204 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net413 net207 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_left_track_13.mux_l1_in_1_ net42 net74 sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk net509
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input39_A chanx_right_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_6.mux_l3_in_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_169_ sb_1__0_.mux_top_track_48.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold68 net512 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold24 net462 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__S sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold35 net466 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 net516 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold57 net536 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold13 net438 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold79 net566 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold340_A sb_1__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_12.mux_l1_in_0_ net41 net105 sb_1__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk
+ net563 net205 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_24.mux_l2_in_0_ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_24.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_6.mux_l2_in_1_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput103 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__buf_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk net382
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.out sky130_fd_sc_hd__clkbuf_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__184__A sb_1__0_.mux_top_track_18.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold302 net353 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold313 sb_1__0_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold357 sb_1__0_.mem_top_track_10.mem_out\[1\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold346 sb_1__0_.mem_top_track_20.mem_out\[0\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold368 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net635
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold324 sb_1__0_.mem_top_track_26.mem_out\[0\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold379 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net646
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold335 sb_1__0_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk net355
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net471
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_24.mux_l1_in_1_ net242 net32 sb_1__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold110 net605 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_right_track_6.mux_l1_in_2_ net16 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_1__0_.mem_right_track_6.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold187 sb_1__0_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold143 net641 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold121 net621 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold198 net297 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold165 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold154 net655 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold132 net629 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold176 net283 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold253_A sb_1__0_.mem_top_track_6.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_0.mux_l1_in_3_ net233 net21 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input69_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold370_A sb_1__0_.mem_right_track_2.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_185_ sb_1__0_.mux_top_track_16.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net208 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk
+ net443 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__0_.mux_left_track_13.mux_l1_in_0_ net66 net78 sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net465
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_168_ sb_1__0_.mux_top_track_50.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_left_track_37.mux_l3_in_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_0.mux_l3_in_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold69 net562 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold14 net430 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 net474 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold58 net548 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold36 net524 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 net460 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chanx_right_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_6.mux_l2_in_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xinput104 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__buf_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_37.mux_l2_in_1_ net217 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input99_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_0.mux_l2_in_1_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_8_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk net402
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold314 sb_1__0_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold347 sb_1__0_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold336 sb_1__0_.mem_top_track_22.mem_out\[0\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold369 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net636
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold358 sb_1__0_.mem_right_track_6.mem_out\[0\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold303 sb_1__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold325 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net592
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_29.mux_l2_in_1__267 VGND VGND VPWR VPWR net267 sb_1__0_.mux_left_track_29.mux_l2_in_1__267/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net575
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net435
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_24.mux_l1_in_0_ net62 net103 sb_1__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__ebufn_8
XFILLER_31_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold144 net647 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold122 net622 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mux_right_track_6.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ net88 sb_1__0_.mem_right_track_6.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold111 net612 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold133 net633 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold100 net602 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 net285 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mux_top_track_36.mux_l2_in_0_ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold199 sb_1__0_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold166 net274 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold155 net657 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold177 sb_1__0_.mem_right_track_20.ccff_tail VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D net499 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_0.mux_l1_in_2_ net24 net51 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_20.mux_l1_in_1__240 VGND VGND VPWR VPWR net240 sb_1__0_.mux_top_track_20.mux_l1_in_1__240/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold363_A sb_1__0_.mem_top_track_0.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__S sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_184_ sb_1__0_.mux_top_track_18.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__S sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input81_A chany_top_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_36.mux_l1_in_1_ net248 net14 sb_1__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_ net261 sb_1__0_.mux_left_track_53.out
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
X_167_ net19 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold26 net490 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 net510 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold15 net446 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold37 net492 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold48 net508 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A chanx_right_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_16.mux_l2_in_1__237 VGND VGND VPWR VPWR net237 sb_1__0_.mux_top_track_16.mux_l2_in_1__237/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net469
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l3_in_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_4.mux_l2_in_1__249 VGND VGND VPWR VPWR net249 sb_1__0_.mux_top_track_4.mux_l2_in_1__249/LO
+ sky130_fd_sc_hd__conb_1
Xinput105 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_37.mux_l2_in_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_0.mux_l2_in_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net513
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold326 sb_1__0_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 sb_1__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold304 net352 VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold359 sb_1__0_.mem_top_track_14.mem_out\[1\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold348 sb_1__0_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net398
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold337 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net604
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_36.mux_l1_in_1__248 VGND VGND VPWR VPWR net248 sb_1__0_.mux_top_track_36.mux_l1_in_1__248/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net533
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_6.mux_l3_in_0__S sb_1__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l2_in_1_ net224 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_6.mux_l1_in_0_ net70 net82 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold167 sb_1__0_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold112 net616 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold145 net644 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold123 net625 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold156 net271 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold101 net598 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold134 net634 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_37.mux_l1_in_1_ net38 net87 sb_1__0_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xhold189 sb_1__0_.mem_top_track_16.mem_out\[0\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold178 net279 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_top_track_0.mux_l1_in_1_ net53 net103 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__ebufn_8
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_183_ sb_1__0_.mux_top_track_20.out VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_12.mux_l1_in_2_ net26 net12 sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_36.mux_l1_in_0_ net44 net105 sb_1__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__S cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_7.mux_l2_in_1__221 VGND VGND VPWR VPWR net221 sb_1__0_.mux_left_track_7.mux_l2_in_1__221/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_top_track_48.mux_l2_in_0_ net254 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__S sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_166_ net20 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_50.mux_l2_in_0_ net255 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_50.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold27 net470 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold38 net530 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold16 net442 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold49 net502 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_24_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold319_A sb_1__0_.mem_right_track_12.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input37_A chanx_right_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net459
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_149_ sb_1__0_.mux_right_track_28.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput106 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_ sb_1__0_.mux_left_track_29.out net9
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__D net479 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold349 sb_1__0_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold305 sb_1__0_.mem_left_track_1.mem_out\[1\] VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold327 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net594
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold338 sb_1__0_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold316 net357 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net401
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold386_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__D net402 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_12.mux_l2_in_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold168 net277 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold113 net615 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold102 net595 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold157 sb_1__0_.mem_top_track_58.mem_out\[0\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold179 sb_1__0_.mem_top_track_18.ccff_tail VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold146 net643 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold135 net631 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold124 net632 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_37.mux_l1_in_0_ net69 net81 sb_1__0_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_0.mux_l1_in_0_ net100 net105 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net207
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_10.mux_l1_in_3__223 VGND VGND VPWR VPWR net223 sb_1__0_.mux_right_track_10.mux_l1_in_3__223/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold349_A sb_1__0_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ sb_1__0_.mux_top_track_22.out VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ net86 sb_1__0_.mem_right_track_12.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input67_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk net499
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__D net539 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_165_ net22 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__S sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 net506 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net496 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold17 net448 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_0__S sb_1__0_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ net9 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_48.mux_l1_in_0_ net10 net103 sb_1__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_6.mux_l2_in_1__A0 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_50.mux_l1_in_0_ net15 net104 sb_1__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold328 sb_1__0_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold306 net348 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold339 sb_1__0_.mem_right_track_4.mem_out\[0\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold317 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net584
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net445
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk net365
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold281_A sb_1__0_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input97_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__S sb_1__0_.mem_top_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold169 sb_1__0_.mem_top_track_4.ccff_tail VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold125 net627 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold158 net272 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold103 net603 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold114 net608 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold147 net646 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold136 net635 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__D net531 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__S sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk net396
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_0__S sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ sb_1__0_.mux_top_track_24.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net409
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l2_in_1__S sb_1__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_12.mux_l1_in_0_ net68 net80 sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk net453
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_42.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout210 net215 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_2
Xsb_1__0_.mux_right_track_36.mux_l3_in_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_164_ sb_1__0_.mux_top_track_58.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net107 net97 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold29 net498 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold18 net454 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__S sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__106__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_147_ net8 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk net531
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk net373
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_21_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.mux_l2_in_1_ net228 net8 sb_1__0_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_ sb_1__0_.mux_left_track_11.out net19
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold157_A sb_1__0_.mem_top_track_58.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input42_A chanx_right_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold329 sb_1__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold307 sb_1__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold318 sb_1__0_.mem_right_track_28.ccff_tail VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net455
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xinput90 chany_top_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 net609 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold126 net617 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold104 net606 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mux_top_track_18.mux_l3_in_0_ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__S sb_1__0_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.out sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold137 net638 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold148 net645 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xhold159 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.out sky130_fd_sc_hd__clkbuf_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net363
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__114__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_180_ sb_1__0_.mux_top_track_26.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk net503
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_18.mux_l2_in_1_ net238 net7 sb_1__0_.mem_top_track_18.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk net553
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_42.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__109__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout211 net215 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_6
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold354_A sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_163_ sb_1__0_.mux_right_track_0.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold19 net452 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk net384
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_5.mux_l3_in_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__122__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_146_ net7 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_1__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net410
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net364
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__S sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0 net35 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.mux_l2_in_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk net501
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_ sb_1__0_.mux_left_track_5.out net22
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_8_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chanx_right_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_21.mux_l3_in_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold308 net345 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA__117__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ net51 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 sb_1__0_.mem_right_track_12.mem_out\[0\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net523
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput91 chany_top_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_1__0_.mux_left_track_5.mux_l2_in_1_ net219 top_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_1__0_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput80 chany_top_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_0__S sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_36.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ net63 sb_1__0_.mem_right_track_36.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_48.mux_l2_in_0__254 VGND VGND VPWR VPWR net254 sb_1__0_.mux_top_track_48.mux_l2_in_0__254/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk net387
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold116 net610 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold149 net648 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 net636 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold105 net604 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold127 net620 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_8_0_prog_clk net439 net209 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_left_track_21.mux_l2_in_1_ net266 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net529
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l3_in_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_13.mux_l2_in_1__265 VGND VGND VPWR VPWR net265 sb_1__0_.mux_left_track_13.mux_l2_in_1__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_18.mux_l2_in_0_ net33 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_18.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__125__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_28.mux_l2_in_1__227 VGND VGND VPWR VPWR net227 sb_1__0_.mux_right_track_28.mux_l2_in_1__227/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__S sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__S sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_20.mux_l2_in_0_ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_21.mux_l1_in_2_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net55 sb_1__0_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xfanout212 net215 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__S sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l2_in_1_ net225 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_162_ sb_1__0_.mux_right_track_2.out VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input65_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk net457
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xinput1 net656 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__S sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_145_ sb_1__0_.mux_right_track_36.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output171_A net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net521
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__0_.mux_top_track_20.mux_l1_in_1_ net240 net5 sb_1__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_33_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk net449
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk net485
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_2.mux_l1_in_2_ net32 net18 sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold309 sb_1__0_.mem_right_track_12.ccff_tail VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkdlybuf4s25_1
X_128_ sb_1__0_.mux_left_track_11.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_5.mux_l2_in_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput92 chany_top_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
Xinput81 chany_top_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput70 chany_top_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout215_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1 net58 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.mux_l1_in_0_ net65 net77 sb_1__0_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk net371
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xhold128 net630 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold106 net601 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold117 net619 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold139 net640 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__S sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_21.mux_l2_in_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold377_A cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input95_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_5.mux_l1_in_1_ net60 net47 sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_21.mux_l1_in_1_ net41 net85 sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xfanout213 net214 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l2_in_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_161_ sb_1__0_.mux_right_track_4.out VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input58_A chanx_right_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__136__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net505
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 net651 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_18.mux_l1_in_0_ net37 net100 sb_1__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_144_ net5 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_14.mux_l2_in_1__236 VGND VGND VPWR VPWR net236 sb_1__0_.mux_top_track_14.mux_l2_in_1__236/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_20.mux_l1_in_0_ net35 net101 sb_1__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_2.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ net90 sb_1__0_.mem_right_track_2.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_32.mux_l2_in_0_ net246 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_127_ sb_1__0_.mux_left_track_13.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout208_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput82 chany_top_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput71 chany_top_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_1.mux_l1_in_3__263 VGND VGND VPWR VPWR net263 sb_1__0_.mux_left_track_1.mux_l1_in_3__263/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chanx_right_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net481
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__144__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 net618 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold129 net624 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold107 net607 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_39_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input88_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_5.mux_l1_in_0_ net92 net75 sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__139__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_0__S sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_21.mux_l1_in_0_ net67 net79 sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xfanout214 net215 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_6
Xfanout203 net208 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_8
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ sb_1__0_.mux_right_track_6.out VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_6.mux_l3_in_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold290 net342 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_45.mux_l3_in_0_ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__152__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input105_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_143_ net4 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input70_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__147__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l1_in_0_ net72 net84 sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_0.mux_l2_in_1__S sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_6.mux_l2_in_1_ net257 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_30 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk net343
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput170 net170 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_ net262 net56 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_45.mux_l2_in_1_ net218 net37 sb_1__0_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_126_ net48 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput72 chany_top_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput83 chany_top_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input33_A chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold108 net611 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_2_ net16 net46 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold119 net626 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkdlybuf4s50_1
X_109_ net59 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_32.mux_l1_in_0_ net26 net56 sb_1__0_.mem_top_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_ net62 net31 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_44.mux_l2_in_0_ net252 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ net350 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__155__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X net108 VGND VGND
+ VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net483
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout204 net208 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_8
Xfanout215 net98 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold291 sb_1__0_.mem_top_track_44.mem_out\[0\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold280 net332 VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__S sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_142_ net32 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input63_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_2.mux_l2_in_1__239 VGND VGND VPWR VPWR net239 sb_1__0_.mux_top_track_2.mux_l2_in_1__239/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_6.mux_l2_in_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net393
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_ net25 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_20.mux_l3_in_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xoutput171 net171 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
Xoutput160 net160 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_45.mux_l2_in_0_ net88 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ net47 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput84 chany_top_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 chany_top_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ net58 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold109 net613 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_1_ net49 net103 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_20.mux_l2_in_1_ net226 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_ net39 net8 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ net403 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout213_A net214 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net429
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_34.mux_l2_in_0__247 VGND VGND VPWR VPWR net247 sb_1__0_.mux_top_track_34.mux_l2_in_0__247/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input93_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_20.mux_l1_in_2_ net25 net11 sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_44.mux_l1_in_0_ net31 net101 sb_1__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout205 net206 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_8
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold281 sb_1__0_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold292 net333 VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold270 net324 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_36_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold240_A net295 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l2_in_1__224 VGND VGND VPWR VPWR net224 sb_1__0_.mux_right_track_12.mux_l2_in_1__224/LO
+ sky130_fd_sc_hd__conb_1
X_141_ sb_1__0_.mux_right_track_44.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input56_A chanx_right_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net569
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_32 sb_1__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput161 net161 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_124_ net46 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__174__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput74 chany_top_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput63 chany_top_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput85 chany_top_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk net573
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_107_ sb_1__0_.mux_left_track_53.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_0_ net100 net105 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__S sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_20.mux_l2_in_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_8_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout206_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_45.mux_l1_in_0_ net70 net82 sb_1__0_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net408 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold320_A sb_1__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__S sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_20.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ net85 sb_1__0_.mem_right_track_20.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout206 net208 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_6
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold271 sb_1__0_.mem_top_track_2.ccff_tail VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold260 net330 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold282 net325 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold293 sb_1__0_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__S sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_140_ net30 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input49_A chanx_right_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_14.mux_l3_in_0_ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_33 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput151 net151 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
XFILLER_28_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__S sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input103_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_123_ sb_1__0_.mux_left_track_21.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l1_in_3_ net263 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput64 chany_top_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 chany_top_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_1
Xinput75 chany_top_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_46.mux_l2_in_0__253 VGND VGND VPWR VPWR net253 sb_1__0_.mux_top_track_46.mux_l2_in_0__253/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_14.mux_l2_in_1_ net236 net9 sb_1__0_.mem_top_track_14.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net415
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_106_ net56 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_ sb_1__0_.mux_left_track_7.out net21
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net487 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold313_A sb_1__0_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_1.mux_l3_in_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_20.mux_l1_in_0_ net67 net79 sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input79_A chany_top_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout207 net208 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_8
Xsb_1__0_.mux_left_track_45.mux_l2_in_1__218 VGND VGND VPWR VPWR net218 sb_1__0_.mux_left_track_45.mux_l2_in_1__218/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_3_0_prog_clk net368
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold261 sb_1__0_.mem_top_track_10.ccff_head VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold283 sb_1__0_.mem_top_track_12.mem_out\[0\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold272 net341 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold250 net313 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold294 net340 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold380_A sb_1__0_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__193__A sb_1__0_.mux_top_track_0.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l2_in_1_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_right_track_44.mux_l1_in_1__230 VGND VGND VPWR VPWR net230 sb_1__0_.mux_right_track_44.mux_l1_in_1__230/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__188__A sb_1__0_.mux_top_track_10.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net376
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_12 net257 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_50.mux_l2_in_0__255 VGND VGND VPWR VPWR net255 sb_1__0_.mux_top_track_50.mux_l2_in_0__255/LO
+ sky130_fd_sc_hd__conb_1
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_28_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__S sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_122_ net43 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input61_A chanx_right_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l1_in_2_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net34 sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 chany_top_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput65 chany_top_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput87 chany_top_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
Xinput98 prog_reset VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ net55 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_14.mux_l2_in_0_ net61 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_14.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk net545
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_ sb_1__0_.mux_left_track_1.out net24
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_0__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout211_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk net425
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout208 net215 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_4
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net374
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold240 net295 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold295 cbx_1__0_.cbx_8__0_.ccff_head VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold262 net331 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold284 net339 VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold273 sb_1__0_.mem_top_track_14.mem_out\[0\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold251 sb_1__0_.mem_right_track_36.ccff_tail VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold373_A sb_1__0_.mem_right_track_10.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input91_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__S sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l2_in_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk net507
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_12.mux_l2_in_1__235 VGND VGND VPWR VPWR net235 sb_1__0_.mux_top_track_12.mux_l2_in_1__235/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk net447
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_13 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_44.mux_l2_in_0_ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_24 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_121_ net42 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input54_A chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_left_track_1.mux_l1_in_1_ net51 net90 sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput77 chany_top_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 chany_top_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput66 chany_top_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput99 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net99 sky130_fd_sc_hd__buf_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__S cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_0__S sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ net44 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_right_track_44.mux_l1_in_1_ net230 net7 sb_1__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_0__S sb_1__0_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net360
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout204_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net479
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_58.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_14.mux_l1_in_0_ net39 net106 sb_1__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_26.mux_l2_in_0_ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_26.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_output123_A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout209 net215 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_8
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk net451
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold263 sb_1__0_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold230 net306 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold296 net336 VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold274 net322 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold241 sb_1__0_.mem_top_track_50.mem_out\[0\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 sb_1__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold252 net311 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input84_A chany_top_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__262 VGND VGND VPWR VPWR net262 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__262/LO
+ sky130_fd_sc_hd__conb_1
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__S cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__S sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_26.mux_l1_in_1_ net243 net30 sb_1__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net392
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output190_A net190 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_197_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_14 net258 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_25 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput121 net121 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput110 net110 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput143 net143 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
XANTENNA_hold329_A sb_1__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_120_ net41 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input47_A chanx_right_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_1.mux_l1_in_0_ net72 net84 sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput89 chany_top_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput78 chany_top_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
Xinput67 chany_top_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_4.mux_l2_in_1__229 VGND VGND VPWR VPWR net229 sb_1__0_.mux_right_track_4.mux_l2_in_1__229/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input101_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__D net425 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_44.mux_l1_in_0_ net64 net76 sb_1__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__259 VGND VGND VPWR VPWR net259 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__259/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net565
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_2.mux_l3_in_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__D net382 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net649 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_2.mux_l2_in_1_ net239 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xhold231 sb_1__0_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold242 net315 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold253 sb_1__0_.mem_top_track_6.ccff_tail VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold220 net309 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 net305 VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold286 net328 VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold275 sb_1__0_.mem_right_track_44.mem_out\[0\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold297 sb_1__0_.mem_top_track_24.ccff_tail VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_28.mux_l2_in_0__244 VGND VGND VPWR VPWR net244 sb_1__0_.mux_top_track_28.mux_l2_in_0__244/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input77_A chany_top_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_26.mux_l1_in_0_ net60 net104 sb_1__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net549
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_2.mux_l1_in_2_ net18 net48 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__S sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_26 net369 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput177 net177 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk net389
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput122 net122 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_40.mux_l2_in_0_ net250 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_1__S sb_1__0_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk net461 net208 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_179_ sb_1__0_.mux_top_track_28.out VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput79 chany_top_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput68 chany_top_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_0__S sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__104__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 net418 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_top_track_32.mux_l2_in_0__246 VGND VGND VPWR VPWR net246 sb_1__0_.mux_top_track_32.mux_l2_in_0__246/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__S sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk net366
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_2.mux_l2_in_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold254 net329 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold265 sb_1__0_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold210 net299 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__S sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold221 sb_1__0_.mem_top_track_16.ccff_tail VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 sb_1__0_.mem_top_track_20.ccff_tail VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold243 sb_1__0_.mem_top_track_18.mem_out\[0\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold232 net296 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold276 net308 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold298 net349 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_53.mux_l3_in_0_ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X cbx_1__0_.cbx_8__0_.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk net361
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold371_A sb_1__0_.mem_right_track_0.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_36.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__112__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_2.mux_l1_in_1_ net52 net104 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_16 chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net385
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_27 chany_top_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0 net41 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
XFILLER_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk net559
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_53.mux_l2_in_1_ net220 net35 sb_1__0_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_19_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_178_ sb_1__0_.mux_top_track_30.out VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput69 chany_top_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold334_A sb_1__0_.mem_top_track_8.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input52_A chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk net491
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_40.mux_l1_in_0_ net3 net99 sb_1__0_.mem_top_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.out sky130_fd_sc_hd__clkbuf_1
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__120__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 net654 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__S sb_1__0_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__115__A sb_1__0_.mux_left_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net406
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xhold255 sb_1__0_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold266 net310 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold222 net321 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold288 net337 VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold233 sb_1__0_.mem_top_track_48.mem_out\[0\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold200 net302 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold244 net326 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold211 sb_1__0_.mem_top_track_50.ccff_tail VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold299 sb_1__0_.mem_top_track_26.ccff_tail VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold277 sb_1__0_.mem_left_track_1.ccff_head VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net551
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_58.mux_l2_in_0__A0 net256 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold364_A sb_1__0_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A chany_top_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_194_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_2.mux_l1_in_0_ net101 net106 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net539
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_28 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_17 chany_top_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput179 net179 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk net495
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_53.mux_l2_in_0_ net89 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
X_177_ sb_1__0_.mux_top_track_32.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_1__0_.mux_right_track_2.mux_l2_in_1__225 VGND VGND VPWR VPWR net225 sb_1__0_.mux_right_track_2.mux_l2_in_1__225/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__S sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_44.mux_l2_in_0__252 VGND VGND VPWR VPWR net252 sb_1__0_.mux_top_track_44.mux_l2_in_0__252/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk net400
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input45_A chanx_right_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__118__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net404
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net208 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__S sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 net422 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_5.mux_l2_in_1__219 VGND VGND VPWR VPWR net219 sb_1__0_.mux_left_track_5.mux_l2_in_1__219/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_10.mux_l3_in_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net517
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xhold201 sb_1__0_.mem_top_track_24.mem_out\[0\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold256 net317 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold223 sb_1__0_.mem_right_track_0.mem_out\[1\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold245 sb_1__0_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold234 net323 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold212 net319 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold267 sb_1__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold278 net334 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold289 sb_1__0_.mem_top_track_46.mem_out\[0\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk net377
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__126__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__S sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net431
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__S sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ sb_1__0_.mux_top_track_0.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_10.mux_l2_in_1_ net234 net12 sb_1__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l1_in_3_ net264 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input75_A chany_top_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 sb_1__0_.mem_left_track_21.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_29 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput125 net125 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
X_176_ sb_1__0_.mux_top_track_34.out VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk net511
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input38_A chanx_right_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net588
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
X_159_ net21 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XANTENNA__134__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_53.mux_l1_in_0_ net71 net83 sb_1__0_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l3_in_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_26.mux_l1_in_1__243 VGND VGND VPWR VPWR net243 sb_1__0_.mux_top_track_26.mux_l1_in_1__243/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 net424 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__129__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0 net62 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_11.mux_l2_in_1_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold235 sb_1__0_.mem_top_track_0.ccff_tail VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold224 net293 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold213 sb_1__0_.mem_right_track_2.ccff_tail VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold202 net290 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold246 net335 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold257 sb_1__0_.mem_top_track_40.mem_out\[0\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold279 sb_1__0_.mem_right_track_10.ccff_tail VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold268 net338 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net390
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__260 VGND VGND VPWR VPWR net260 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__260/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__142__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__ebufn_8
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_192_ sb_1__0_.mux_top_track_2.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_10.mux_l2_in_1__234 VGND VGND VPWR VPWR net234 sb_1__0_.mux_top_track_10.mux_l2_in_1__234/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_10.mux_l2_in_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l1_in_2_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net58 sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input68_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput115 net115 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_175_ sb_1__0_.mux_top_track_36.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_10.mux_l1_in_1_ net40 net42 sb_1__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net489
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_158_ sb_1__0_.mux_right_track_10.out VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__150__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input50_A chanx_right_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 net426 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_7.mux_l3_in_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net537
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold282_A net325 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input98_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_11.mux_l2_in_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xhold203 sb_1__0_.mem_left_track_53.mem_out\[0\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold236 net316 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold214 net300 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold225 sb_1__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold258 net303 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold269 sb_1__0_.mem_top_track_30.mem_out\[0\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold247 sb_1__0_.mem_top_track_28.mem_out\[0\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net473
+ net210 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_7.mux_l2_in_1_ net221 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__S sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1 net56 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ sb_1__0_.mux_top_track_4.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_left_track_11.mux_l1_in_1_ net43 net63 sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mux_right_track_4.mux_l3_in_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_3_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_7.mux_l1_in_2_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ top_width_0_height_0_subtile_0__pin_inpad_0_ sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__ebufn_8
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input80_A chany_top_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ net362 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_174_ net106 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__148__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0 sb_1__0_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_10.mux_l1_in_0_ net102 net99 sb_1__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_0__S sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_22.mux_l2_in_0_ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_22.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_157_ sb_1__0_.mux_right_track_12.out VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_4.mux_l2_in_1_ net229 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input43_A chanx_right_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold7 net432 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net583
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_22.mux_l1_in_1_ net241 net4 sb_1__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_4.mux_l1_in_2_ net30 net17 sb_1__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__156__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold204 net294 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold237 sb_1__0_.mem_top_track_14.ccff_tail VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold226 net304 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold259 sb_1__0_.mem_top_track_32.mem_out\[0\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold248 net318 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold215 sb_1__0_.mem_top_track_34.mem_out\[0\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_7.mux_l2_in_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ sb_1__0_.mux_top_track_6.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net397
+ net208 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_11.mux_l1_in_0_ net65 net77 sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_8.mux_l2_in_1__258 VGND VGND VPWR VPWR net258 sb_1__0_.mux_top_track_8.mux_l2_in_1__258/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_58.mux_l2_in_0__256 VGND VGND VPWR VPWR net256 sb_1__0_.mux_top_track_58.mux_l2_in_0__256/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_0__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput117 net117 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_52.mux_l2_in_0_ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_7.mux_l1_in_1_ net59 net46 sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_173_ sb_1__0_.mux_top_track_40.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ net391 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_right_track_0.mux_l2_in_1__222 VGND VGND VPWR VPWR net222 sb_1__0_.mux_right_track_0.mux_l2_in_1__222/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_156_ net18 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_52.mux_l1_in_1_ net231 net5 sb_1__0_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_4.mux_l2_in_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__159__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chanx_right_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 net428 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_15_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_139_ net29 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_30.mux_l2_in_0__245 VGND VGND VPWR VPWR net245 sb_1__0_.mux_top_track_30.mux_l2_in_0__245/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_22.mux_l1_in_0_ net34 net102 sb_1__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_4.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ net89 sb_1__0_.mem_right_track_4.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_3.mux_l2_in_1__216 VGND VGND VPWR VPWR net216 sb_1__0_.mux_left_track_3.mux_l2_in_1__216/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_top_track_34.mux_l2_in_0_ net247 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold238 net312 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold227 sb_1__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold205 sb_1__0_.mem_right_track_4.ccff_tail VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold249 sb_1__0_.mem_right_track_10.ccff_head VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold216 net298 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_6.mux_l1_in_3__232 VGND VGND VPWR VPWR net232 sb_1__0_.mux_right_track_6.mux_l1_in_3__232/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_0__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__S sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__D net435 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_3_ net223 net28 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net535
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net207 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput107 net107 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XFILLER_9_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput118 net118 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
XFILLER_36_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_ net259 net59 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_7.mux_l1_in_0_ net64 net76 sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_0__S sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net414 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ sb_1__0_.mux_top_track_42.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input66_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__180__A sb_1__0_.mux_top_track_26.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_155_ net17 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_52.mux_l1_in_0_ net92 net75 sb_1__0_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_10.mux_l3_in_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_ sb_1__0_.mux_left_track_37.out net5
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_8.mux_l3_in_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA__175__A sb_1__0_.mux_top_track_36.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold9 net440 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_138_ net28 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_0__S sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_10.mux_l2_in_1_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_4.mux_l1_in_0_ net71 net83 sb_1__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_8.mux_l2_in_1_ net258 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_8.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold206 net301 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold217 sb_1__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold239 sb_1__0_.mem_left_track_29.mem_out\[1\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold228 net307 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk net379
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold378_A sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input96_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A0 sb_1__0_.mux_left_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_2_ net13 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_right_track_10.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_34.mux_l1_in_0_ net25 net55 sb_1__0_.mem_top_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_8.mux_l1_in_2_ net13 net43 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__S sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput119 net119 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mux_top_track_46.mux_l2_in_0_ net253 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput108 net108 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk
+ net427 net204 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ sb_1__0_.mux_top_track_44.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk net367
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_42.mux_l2_in_0__251 VGND VGND VPWR VPWR net251 sb_1__0_.mux_top_track_42.mux_l2_in_0__251/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__S sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold360_A sb_1__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_154_ net16 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_53.mux_l2_in_1__220 VGND VGND VPWR VPWR net220 sb_1__0_.mux_left_track_53.mux_l2_in_1__220/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net399
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_137_ sb_1__0_.mux_right_track_52.out VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout209_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold323_A sb_1__0_.mem_right_track_20.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_10.mux_l2_in_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input41_A chanx_right_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_8.mux_l2_in_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xhold229 sb_1__0_.mem_top_track_12.ccff_tail VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold207 sb_1__0_.mem_left_track_1.ccff_tail VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold218 net320 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net383
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input89_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_2_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold90 net582 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ net87 sb_1__0_.mem_right_track_10.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_8.mux_l1_in_1_ net45 net104 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput109 net109 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.out sky130_fd_sc_hd__clkbuf_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_170_ sb_1__0_.mux_top_track_46.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold390 net1 VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_33_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__189__A sb_1__0_.mux_top_track_8.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net359
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__S sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input106_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_46.mux_l1_in_0_ net6 net102 sb_1__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_15_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ sb_1__0_.mux_right_track_20.out VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input71_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_ sb_1__0_.mux_left_track_13.out net18
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_58.mux_l2_in_0_ net256 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_24.mux_l1_in_1__242 VGND VGND VPWR VPWR net242 sb_1__0_.mux_top_track_24.mux_l1_in_1__242/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net370
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net561
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_136_ net26 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input34_A chanx_right_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold208 net314 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkdlybuf4s25_1
X_119_ sb_1__0_.mux_left_track_29.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold219 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__D net549 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk net475
+ net205 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk net433 net208 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold91 net594 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold80 net578 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_0_ net69 net81 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_8.mux_l1_in_0_ net101 net106 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__S sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net206 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold380 sb_1__0_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net577
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_152_ net13 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input64_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_ sb_1__0_.mux_left_track_7.out net21
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__S cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__S sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk net555
+ net211 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net215 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_135_ net25 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__S sb_1__0_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_21.mux_l2_in_1__A0 net266 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold211_A sb_1__0_.mem_top_track_50.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_58.mux_l1_in_0_ net23 net54 sb_1__0_.mem_top_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_16.mux_l3_in_0_ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_118_ net39 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xhold209 sb_1__0_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold70 net554 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold81 net572 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold92 net590 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net515
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_37.mux_l2_in_1__217 VGND VGND VPWR VPWR net217 sb_1__0_.mux_left_track_37.mux_l2_in_1__217/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_16.mux_l2_in_1_ net237 net8 sb_1__0_.mem_top_track_16.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_10_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__D net513 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input94_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk net395
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__S cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 sb_1__0_.mem_right_track_2.mem_out\[0\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold381 ccff_head_1 VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_3.mux_l3_in_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_17_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_151_ net12 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ sb_1__0_.mux_left_track_1.out net24
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input57_A chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_3.mux_l2_in_1_ net216 top_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_1__0_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_134_ net14 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ net38 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout207_A net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_0.mux_l3_in_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold60 net580 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_output126_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold71 net534 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold93 net591 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold82 net564 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net567
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 net235 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_16.mux_l2_in_0_ net57 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_16.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_6.mux_l2_in_1__257 VGND VGND VPWR VPWR net257 sb_1__0_.mux_top_track_6.mux_l2_in_1__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_0.mux_l2_in_1_ net222 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_0.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net411
+ net212 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk net525
+ net204 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_6_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold371 sb_1__0_.mem_right_track_0.mem_out\[0\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold360 sb_1__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold382 net416 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_21.mux_l2_in_1__266 VGND VGND VPWR VPWR net266 sb_1__0_.mux_left_track_21.mux_l2_in_1__266/LO
+ sky130_fd_sc_hd__conb_1
X_150_ net11 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold190 net287 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mux_right_track_0.mux_l1_in_2_ net4 net21 sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l2_in_0__S sb_1__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_right_track_36.mux_l2_in_1__228 VGND VGND VPWR VPWR net228 sb_1__0_.mux_right_track_36.mux_l2_in_1__228/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_hold10_A net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold351_A sb_1__0_.mem_top_track_4.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input104_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk net369
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk net380
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_133_ sb_1__0_.mux_left_track_1.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_left_track_3.mux_l2_in_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__110__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold58_A net548 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__S sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ net37 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XANTENNA__105__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net207
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_29.mux_l3_in_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_3.mux_l1_in_1_ net62 net48 sb_1__0_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold50 net522 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold72 net550 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold94 net597 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold61 net552 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold83 net584 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_3 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__S sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l2_in_1_ net267 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net214 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_0.mux_l2_in_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net419
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net441
+ net203 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 sb_1__0_.mem_left_track_37.mem_out\[0\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold372 sb_1__0_.mem_top_track_2.mem_out\[0\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold383 net268 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_hold381_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold361 sb_1__0_.mem_right_track_28.mem_out\[1\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net381
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__113__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_16.mux_l1_in_0_ net38 net99 sb_1__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_29.mux_l1_in_2_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net44 sb_1__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_28.mux_l2_in_0_ net244 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 net282 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_0.mux_l1_in_1_ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold191 sb_1__0_.mem_top_track_22.ccff_tail VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net543
+ net209 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk net386
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_30.mux_l2_in_0_ net245 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__108__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net378
+ net213 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net388
+ net206 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_132_ sb_1__0_.mux_left_track_3.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input62_A chanx_right_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk net557
+ net207 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_29_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_115_ sb_1__0_.mux_left_track_37.out VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__121__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_3.mux_l1_in_0_ net91 net73 sb_1__0_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk net477
+ net214 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold307_A sb_1__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold40 net494 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold62 net520 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold84 net576 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold51 net514 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold73 net560 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold95 net592 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__116__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout212_A net215 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l2_in_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_4.mux_l3_in_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

