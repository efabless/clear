* NGSPICE file created from tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

.subckt tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0] chanx_right_in_0[10]
+ chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13] chanx_right_in_0[14]
+ chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17] chanx_right_in_0[18]
+ chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20] chanx_right_in_0[21]
+ chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24] chanx_right_in_0[25]
+ chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28] chanx_right_in_0[29]
+ chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4] chanx_right_in_0[5]
+ chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8] chanx_right_in_0[9]
+ chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11] chanx_right_out_0[12]
+ chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15] chanx_right_out_0[16]
+ chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19] chanx_right_out_0[1]
+ chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22] chanx_right_out_0[23]
+ chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26] chanx_right_out_0[27]
+ chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2] chanx_right_out_0[3]
+ chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6] chanx_right_out_0[7]
+ chanx_right_out_0[8] chanx_right_out_0[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] clk0 prog_clk prog_reset reset right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ top_width_0_height_0_subtile_0__pin_O_0_
+ top_width_0_height_0_subtile_0__pin_O_1_ top_width_0_height_0_subtile_0__pin_O_2_
+ top_width_0_height_0_subtile_0__pin_O_3_ top_width_0_height_0_subtile_0__pin_O_4_
+ top_width_0_height_0_subtile_0__pin_O_5_ top_width_0_height_0_subtile_0__pin_O_6_
+ top_width_0_height_0_subtile_0__pin_O_7_ top_width_0_height_0_subtile_0__pin_cin_0_
+ top_width_0_height_0_subtile_0__pin_reg_in_0_
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_1__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_37.mux_l1_in_1_ net68 net38 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_53_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_3__S sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input127_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3_ net306 net116 cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3__411 VGND VGND VPWR VPWR net411 cbx_1__1_.mux_top_ipin_14.mux_l2_in_3__411/LO
+ sky130_fd_sc_hd__conb_1
X_363_ net81 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input92_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_294_ net11 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_1__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_28.mux_l2_in_3__388 VGND VGND VPWR VPWR net388 sb_1__1_.mux_right_track_28.mux_l2_in_3__388/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_1__A0 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_0__S sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l4_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l2_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_91_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_2_ net14 net35 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_13.ccff_tail net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__1_.mem_left_track_3.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_346_ net92 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_277_ sb_1__1_.mux_left_track_1.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net429 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_3__A1 sb_1__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_0.mux_l2_in_3_ net394 net4 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_52_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_28.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput253 net253 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput242 net242 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput231 net231 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput264 net264 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput275 net275 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__328
+ VGND VGND VPWR VPWR net328 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__328/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net441 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l3_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_1_ net65 net130 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input55_A chanx_right_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_3.mux_l1_in_1_ net48 net93 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ net107 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_3.mux_l4_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__buf_4
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_2__A0 sb_1__1_.mux_left_track_21.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_3__S sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3__408 VGND VGND VPWR VPWR net408 cbx_1__1_.mux_top_ipin_11.mux_l2_in_3__408/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3__310 VGND VGND VPWR VPWR net310 cby_1__1_.mux_right_ipin_7.mux_l2_in_3__310/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_0__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3__413 VGND VGND VPWR VPWR net413 cbx_1__1_.mux_top_ipin_2.mux_l2_in_3__413/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_2__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA__312__A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net143 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l2_in_2_ net13 sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3_ net311 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_2__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_2__S sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l4_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold41 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR
+ net454 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold30 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X VGND VGND VPWR VPWR
+ net443 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold63 net421 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold52 sb_1__1_.mem_left_track_37.ccff_tail VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_0__S sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_2__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_1_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_1__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__351
+ VGND VGND VPWR VPWR net351 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__351/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_28.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_1__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_2.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput120 chany_top_in_0[7] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
XFILLER_76_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput131 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xinput142 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_3__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_0__S sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_3_ net75 net132 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_2__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_2__S cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l1_in_0_ net98 net110 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_4__A0 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.mux_l3_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_2_ net85 sb_1__1_.mux_bottom_track_37.out cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_26_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_362_ sb_1__1_.mux_top_track_10.out VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3__307 VGND VGND VPWR VPWR net307 cby_1__1_.mux_right_ipin_4.mux_l2_in_3__307/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_293_ sb_1__1_.mux_right_track_28.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input85_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_2__S sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_1__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l4_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_1_ net4 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_52_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_0__S sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__320__A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_28.mux_l1_in_1_ net44 net61 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_1.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_88_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net353 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_345_ sb_1__1_.mux_top_track_44.out VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
X_276_ sb_1__1_.mux_left_track_3.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_24_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_2_ net21 net24 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__1_.mem_top_track_28.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__354
+ VGND VGND VPWR VPWR net354 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__354/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__315__A sb_1__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput210 net210 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput243 net243 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput221 net221 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
Xoutput254 net254 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput265 net265 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput276 net276 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l3_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_52.mux_l1_in_0_ net117 net95 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net332 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_3__S sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_2_ net41 net10 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input48_A chanx_right_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.out sky130_fd_sc_hd__buf_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_0__S sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_1__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_328_ net106 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
X_259_ sb_1__1_.mux_left_track_37.out VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input102_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_0__S sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_3__S sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_3__A0 sb_1__1_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_0__A0 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l2_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold20 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold31 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X VGND VGND VPWR VPWR
+ net444 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold64 sc_in VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold53 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ net455 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_2__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output271_A net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_20.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net346 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__mux2_4
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA__323__A sb_1__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__320
+ VGND VGND VPWR VPWR net320 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__320/LO
+ sky130_fd_sc_hd__conb_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_2__A0 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_1__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 chany_top_in_0[25] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_2__S sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput121 chany_top_in_0[8] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xinput143 net433 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_42_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l1_in_2_ net130 net128 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__318__A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_4__A1 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.mux_l3_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l2_in_3__A1 sb_1__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_1_ net65 cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_361_ sb_1__1_.mux_top_track_12.out VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_21.mux_l2_in_3_ net375 net285 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
X_292_ net9 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input78_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[2\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_2__S sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_3__A0 sb_1__1_.mux_left_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l1_in_0_ net39 net135 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_0__S sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input132_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ net90 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_1__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_275_ sb_1__1_.mux_left_track_5.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_3__S sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] net287 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_37.mux_l2_in_1__378 VGND VGND VPWR VPWR net378 sb_1__1_.mux_left_track_37.mux_l2_in_1__378/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_1__S sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3__292 VGND VGND VPWR VPWR net292 cbx_1__1_.mux_top_ipin_5.mux_l2_in_3__292/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_91_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_top_track_28.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xoutput200 net200 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput244 net244 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput255 net255 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput266 net266 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__331__A sb_1__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput277 net277 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_4__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_2.mux_l2_in_3_ net386 net32 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_327_ sb_1__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_258_ net35 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_0__A0 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_3__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_21.mux_l4_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA__326__A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_0.mux_l1_in_2_ net34 net51 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_0__S sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__332
+ VGND VGND VPWR VPWR net332 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__332/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_84_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l2_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_37_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold21 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold10 net425 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold32 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ net445 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold43 chany_bottom_in[16] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_2__A0 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_2__A0 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_21.mux_l3_in_1_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l4_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__340
+ VGND VGND VPWR VPWR net340 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__340/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 chany_top_in_0[16] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 chany_top_in_0[26] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_4
XFILLER_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput122 chany_top_in_0[9] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_4
Xinput133 net426 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 net428 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_2__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l1_in_1_ net126 net118 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_0__S sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net342 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_2__S sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__334__A sb_1__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_45_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_0__S sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_360_ net78 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_21.mux_l2_in_2_ net279 net85 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_291_ net8 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3_ net290 net56 cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_2.mux_l3_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__329__A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input125_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_343_ net89 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_1__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ sb_1__1_.mux_left_track_7.out VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input90_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_3_ net396 net26 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[0\] net287 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_76_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput201 net201 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput234 net234 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput256 net256 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput245 net245 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput267 net267 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput278 net278 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_2_ net18 net91 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net350 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_2.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__344
+ VGND VGND VPWR VPWR net344 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__344/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_326_ net103 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_257_ net34 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_0__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_bottom_track_3.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_3__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA__342__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_0__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_0.mux_l1_in_1_ net53 net139 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__252__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input53_A chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_61_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_3__S sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_309_ net115 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_2__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_0__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_0__S sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__337__A sb_1__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.mux_l4_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3_ net295 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold22 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_3__S sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold11 net124 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_12
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold44 cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ net457 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_2__A1 net278 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_2__A1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_1__S cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_21.mux_l3_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_74_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_3__A0 sb_1__1_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3_ net365 net14 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_0__A0 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput101 chany_top_in_0[17] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput112 chany_top_in_0[27] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput134 net431 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_6
Xinput123 net417 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_1_0__f_clk0_A clknet_0_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net328 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__mux2_4
XFILLER_8_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_0_ net103 net110 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_12.mux_l3_in_1_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__350__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ net7 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_1_ net71 sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_2_ net25 sb_1__1_.mux_left_track_37.out cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_1__A0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__260__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_0__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_11.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[0\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l3_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_2__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__333
+ VGND VGND VPWR VPWR net333 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__333/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_8.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__356
+ VGND VGND VPWR VPWR net356 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__356/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input118_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_342_ net88 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_273_ net51 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XANTENNA__255__A sb_1__1_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input83_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_2_ net10 net12 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ net470 net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_29.mux_l4_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput213 net213 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput235 net235 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput246 net246 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput268 net268 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput257 net257 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_3__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput279 net279 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_21.mux_l1_in_2_ net75 net55 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_1__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_2.mux_l2_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_12.mux_l2_in_3__385 VGND VGND VPWR VPWR net385 sb_1__1_.mux_right_track_12.mux_l2_in_3__385/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_51_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_2.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ net102 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_256_ net62 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_1__S sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_0.mux_l1_in_0_ net136 net141 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_1_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input46_A chanx_right_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_1__S sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_11.mux_l2_in_3__373 VGND VGND VPWR VPWR net373 sb_1__1_.mux_left_track_11.mux_l2_in_3__373/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ net104 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_2__A1 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.mux_l1_in_2_ net132 net129 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3__303 VGND VGND VPWR VPWR net303 cby_1__1_.mux_right_ipin_14.mux_l2_in_3__303/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_0__A0 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold23 chany_bottom_in[0] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold12 reset VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 chanx_left_in[12] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold34 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input100_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__263__A sb_1__1_.mux_left_track_29.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__348__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_2_ net31 net9 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_1__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_0__A1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput102 chany_top_in_0[18] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
Xinput135 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput113 chany_top_in_0[28] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput124 net423 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_6
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_2__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__258__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l3_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_0_prog_clk net466 net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3__365 VGND VGND VPWR VPWR net365 sb_1__1_.mux_bottom_track_29.mux_l2_in_3__365/LO
+ sky130_fd_sc_hd__conb_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_21.mux_l2_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_1_ net5 cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_11.ccff_head
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net357 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_tail net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_1__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3__298 VGND VGND VPWR VPWR net298 cby_1__1_.mux_right_ipin_1.mux_l2_in_3__298/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_41_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_1__A0 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_2__S sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_1__S sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_341_ sb_1__1_.mux_top_track_52.out VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ sb_1__1_.mux_left_track_11.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_1_ net86 sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__271__A sb_1__1_.mux_left_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input76_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput203 net203 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput214 net214 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput258 net258 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput247 net247 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput236 net236 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput269 net269 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_left_track_21.mux_l1_in_1_ net41 net115 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__356__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net323 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_0__S sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_2.mux_l2_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_2.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input130_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__266__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ net101 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_255_ sb_1__1_.mux_left_track_45.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3_ net299 net115 cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_12.mux_l1_in_2_ net72 net56 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_3__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_52.mux_l2_in_1__392 VGND VGND VPWR VPWR net392 sb_1__1_.mux_right_track_52.mux_l2_in_1__392/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_2__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chanx_right_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_307_ sb_1__1_.mux_right_track_0.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_1__A0 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l1_in_1_ net126 net122 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold13 net477 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold35 chany_bottom_in[4] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 chanx_left_in[13] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold24 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X VGND VGND VPWR VPWR
+ net437 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold57 sb_1__1_.mem_bottom_track_37.ccff_tail VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_2.mux_l2_in_3__397 VGND VGND VPWR VPWR net397 sb_1__1_.mux_top_track_2.mux_l2_in_3__397/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_2__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_1_ net269 net44 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_1__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput103 chany_top_in_0[19] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xinput136 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput114 chany_top_in_0[29] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput125 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net125 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__274__A sb_1__1_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_10.mux_l4_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__359__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_3__S sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__329
+ VGND VGND VPWR VPWR net329 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__329/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3__305 VGND VGND VPWR VPWR net305 cby_1__1_.mux_right_ipin_2.mux_l2_in_3__305/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__269__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__322
+ VGND VGND VPWR VPWR net322 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__322/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3_ net304 net122 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_1__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_2__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_340_ net86 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ sb_1__1_.mux_left_track_13.out VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input69_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xoutput204 net204 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput248 net248 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput259 net259 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput237 net237 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_21.mux_l1_in_0_ net101 net105 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_36.mux_l2_in_1__400 VGND VGND VPWR VPWR net400 sb_1__1_.mux_top_track_36.mux_l2_in_1__400/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_2__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_2__S sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_55_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_3__A1 net285 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_0.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_323_ sb_1__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
X_254_ net60 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__282__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3_ net411 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__D cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.mux_l3_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l1_in_1_ net40 net42 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_0__S sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_15.mux_l4_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.ccff_tail VGND
+ VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_74_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__277__A sb_1__1_.mux_left_track_1.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_1__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_306_ sb_1__1_.mux_right_track_2.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_1__A1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.mux_l1_in_0_ net108 net114 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__341
+ VGND VGND VPWR VPWR net341 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__341/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_1__S sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_2__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold14 net133 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold47 cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR net460
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xhold25 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X VGND VGND VPWR VPWR
+ net438 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X VGND VGND VPWR VPWR
+ net449 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold58 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_1__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3__369 VGND VGND VPWR VPWR net369 sb_1__1_.mux_bottom_track_5.mux_l2_in_3__369/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_left_track_45.mux_l2_in_1_ net379 sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_1__A0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A chanx_right_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_2__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_2__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_21_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_14.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_1_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput104 chany_top_in_0[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
Xinput115 chany_top_in_0[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput126 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net126 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput137 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net137 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_2__S sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__314
+ VGND VGND VPWR VPWR net314 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__314/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__290__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_3__A0 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_load_slew289_A net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_45.mux_l1_in_2_ net282 net91 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l2_in_3__A1 sb_1__1_.mux_left_track_53.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_1_ net39 net52 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_94_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_2_ net91 net99 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net143 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net339 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__mux2_4
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_3__S sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_270_ net48 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_3__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3__290 VGND VGND VPWR VPWR net290 cbx_1__1_.mux_top_ipin_3.mux_l2_in_3__290/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_0.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput216 net216 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput205 net205 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput249 net249 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput227 net227 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput238 net238 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_2.mux_l2_in_3__386 VGND VGND VPWR VPWR net386 sb_1__1_.mux_right_track_2.mux_l2_in_3__386/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_2__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3_ net307 net115 cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input116_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__336
+ VGND VGND VPWR VPWR net336 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__336/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__315
+ VGND VGND VPWR VPWR net315 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__315/LO
+ sky130_fd_sc_hd__conb_1
X_322_ net99 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
X_253_ net59 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input81_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_12.mux_l1_in_0_ net139 net141 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_3__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_10.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_1__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net359 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_305_ sb_1__1_.mux_right_track_4.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output285_A net285 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_36.mux_l3_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_1__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold15 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold26 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ net439 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xhold37 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X VGND VGND VPWR VPWR
+ net450 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold48 chany_bottom_in[12] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__326
+ VGND VGND VPWR VPWR net326 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__326/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_0__S sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.mux_l2_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_1__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A chanx_right_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__288__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l4_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_3__A1 sb_1__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net313 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l2_in_2__A0 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput105 chany_top_in_0[20] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xinput116 chany_top_in_0[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput127 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput138 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_3__A1 net270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_36.mux_l2_in_1_ net400 sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_94_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3_ net312 net119 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk cby_1__1_.mem_right_ipin_3.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_2__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_45.mux_l1_in_1_ net67 net37 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_36.mux_l2_in_1__389 VGND VGND VPWR VPWR net389 sb_1__1_.mux_right_track_36.mux_l2_in_1__389/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_0_ net104 net99 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_11.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[0\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_36.mux_l1_in_2_ net8 net20 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_3_ net404 net29 sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 net427 net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_13.ccff_tail
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XANTENNA__296__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_1__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput217 net217 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput206 net206 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput239 net239 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput228 net228 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold15_A top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_3__S sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_3__A1 net280 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input109_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_321_ net98 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
X_252_ net58 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l4_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_input74_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_40_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__338
+ VGND VGND VPWR VPWR net338 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__338/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_6.mux_l1_in_4_ net16 net89 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_3__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_304_ sb_1__1_.mux_right_track_6.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output278_A net278 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_7_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l4_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_2__S sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold16 net144 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_6.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xhold27 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold38 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X VGND VGND VPWR VPWR
+ net451 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold49 cby_1__1_.mem_right_ipin_4.ccff_tail VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_1_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_71_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input37_A chanx_right_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_14.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_3__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_1__S sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput106 chany_top_in_0[21] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
Xinput117 chany_top_in_0[4] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput128 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net128 sky130_fd_sc_hd__clkbuf_2
Xinput139 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_1__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_0__A0 sb_1__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_36.mux_l2_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__299__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l3_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_0.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_0__S sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_28.mux_l2_in_3_ net388 net14 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_2__S sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_2_ net88 net99 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold45_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_2__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.mux_l1_in_0_ net97 net112 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_4__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input139_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_0__S sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_0__S sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_2__A0 sb_1__1_.mux_left_track_13.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_2__S sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_29.ccff_tail net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_2__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_0__A0 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3_ net363 net26 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk cbx_1__1_.mem_top_ipin_0.ccff_tail
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_36.mux_l1_in_1_ net68 net57 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_2_ net31 sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_0__S sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_30_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net321 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__mux2_2
Xoutput207 net207 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput229 net229 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net348 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_2__A0 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_28.mux_l4_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_320_ net97 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_2__A0 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_251_ sb_1__1_.mux_left_track_53.out VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input67_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l1_in_3_ net76 net59 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input121_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ net21 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_2__A0 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_4__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_bottom_track_13.mux_l4_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_3__S sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_21.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_1__A0 net272 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3__301 VGND VGND VPWR VPWR net301 cby_1__1_.mux_right_ipin_12.mux_l2_in_3__301/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l3_in_1_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xhold17 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold28 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold39 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_2__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l2_in_3__394 VGND VGND VPWR VPWR net394 sb_1__1_.mux_top_track_0.mux_l2_in_3__394/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_3__S sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_3__S sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__A0 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_53.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_65_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net331 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput107 chany_top_in_0[22] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput118 chany_top_in_0[5] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xinput129 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_1__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_1__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_1_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_3__S sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.ccff_tail
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l3_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_0.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_2_ net9 net74 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_15_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net447 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_top_track_20.mux_l2_in_3__398 VGND VGND VPWR VPWR net398 sb_1__1_.mux_top_track_20.mux_l2_in_3__398/LO
+ sky130_fd_sc_hd__conb_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xload_slew286 net415 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input97_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_load_slew287_A net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_3__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_2_ net10 net12 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_85_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_3__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_2__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_36.mux_l1_in_0_ net38 net136 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_2__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput208 net208 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3__363 VGND VGND VPWR VPWR net363 sb_1__1_.mux_bottom_track_13.mux_l2_in_3__363/LO
+ sky130_fd_sc_hd__conb_1
Xoutput219 net219 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_31_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_6.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_2__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_10.mux_l2_in_3__384 VGND VGND VPWR VPWR net384 sb_1__1_.mux_right_track_10.mux_l2_in_3__384/LO
+ sky130_fd_sc_hd__conb_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3_ net291 net55 cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_86_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_2__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_2__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ net56 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_2__S sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold20_A top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3_ net369 net30 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__358
+ VGND VGND VPWR VPWR net358 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__358/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l1_in_2_ net46 net49 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input114_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3__405 VGND VGND VPWR VPWR net405 cbx_1__1_.mux_top_ipin_0.mux_l2_in_3__405/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_2__S sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_302_ sb_1__1_.mux_right_track_10.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_4__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_6.ccff_tail
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_21.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_5.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_1__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l3_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xhold18 test_enable VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold29 chanx_left_in[1] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3__366 VGND VGND VPWR VPWR net366 sb_1__1_.mux_bottom_track_3.mux_l2_in_3__366/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output283_A net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__A1 net279 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_53.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCD
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput108 chany_top_in_0[23] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
Xinput119 chany_top_in_0[6] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_prog_clk_A clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l4_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_79_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input42_A chanx_right_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_0.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_2__A0 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_1_ net69 net82 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_1__A0 net270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew287 net288 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3_ net296 net59 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 chany_bottom_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[2\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_2__S sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_3__A1 net285 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_12_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_0__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_1_ net273 sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_85_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_1__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_2__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_1_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l2_in_3_ net398 net25 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 net209 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_2__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_0__S sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_84_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_0.mux_l2_in_3__383 VGND VGND VPWR VPWR net383 sb_1__1_.mux_right_track_0.mux_l2_in_3__383/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_6.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_77_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_9.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_0__S sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_2_ net275 net56 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1__370 VGND VGND VPWR VPWR net370 sb_1__1_.mux_bottom_track_53.mux_l2_in_1__370/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_2_ net17 net20 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l1_in_1_ net139 net137 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__359
+ VGND VGND VPWR VPWR net359 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__359/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_1__S sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input107_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ sb_1__1_.mux_right_track_12.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input72_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_left_track_21.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_73_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_5.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xhold19 net134 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_12
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_20.mux_l4_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net329 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_3__A0 sb_1__1_.mux_left_track_29.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_1__A0 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l2_in_3_ net380 net283 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_21_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output276_A net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_45.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net349 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput109 chany_top_in_0[24] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_2__S sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input35_A chanx_right_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk net422
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_2__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_28.mux_l2_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_7.mux_l2_in_3__382 VGND VGND VPWR VPWR net382 sb_1__1_.mux_left_track_7.mux_l2_in_3__382/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_3__S sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_2__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_20.mux_l3_in_1_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xload_slew288 net415 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__buf_12
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_2_ net28 net39 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_3__A0 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net320 net434 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xinput91 chany_bottom_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput80 chany_bottom_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[1\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_1__S sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_0__A1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_0__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_3__S sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold43_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__310__A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l4_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_0__S sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_4__S sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_28.mux_l1_in_1_ net127 net104 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input137_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_20.mux_l2_in_2_ net11 net15 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_2__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_1__S sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_6.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net358 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__mux2_2
XFILLER_10_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_3__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_1_ net42 net49 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_0__A0 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_1_ net272 sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l3_in_1_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_95_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_6.mux_l1_in_0_ net135 net141 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_0__S cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_91_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_1__A0 net272 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_300_ net18 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input65_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_0__S sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net440 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_5.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 net474 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_10_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3__361 VGND VGND VPWR VPWR net361 sb_1__1_.mux_bottom_track_1.mux_l2_in_3__361/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__323
+ VGND VGND VPWR VPWR net323 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__323/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3__295 VGND VGND VPWR VPWR net295 cbx_1__1_.mux_top_ipin_8.mux_l2_in_3__295/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_2_ net269 net60 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l2_in_2_ net280 net90 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_7_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output269_A net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_61_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3_ net300 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__313__A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput190 net190 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
XFILLER_94_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_1__S sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l3_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xload_slew289 net415 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_16
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__308__A net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_3__A1 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput70 net456 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xinput81 chany_bottom_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[0\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput92 chany_bottom_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_69_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3_ net407 net55 cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__331
+ VGND VGND VPWR VPWR net331 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__331/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_1__S sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_3__S cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ net445 VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_28.mux_l1_in_0_ net99 net100 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCD
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l4_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input95_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_0__A0 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_20.mux_l2_in_1_ net85 sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_1__S sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__321__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_10.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_3__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_0__S sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk net467 net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net318 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_0_ net116 net102 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_70_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_2__A0 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_5.mux_l3_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__318
+ VGND VGND VPWR VPWR net318 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__318/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_36_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__316__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_1_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_86_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_20.mux_l1_in_2_ net71 net55 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_37.mux_l3_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_4__S sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chanx_right_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_1__S sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_60_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_359_ net77 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net146 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_0__S sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput2 net476 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3_ net412 net62 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_input112_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_1_ net36 net47 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_1_ net77 sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_1__A0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_1__S sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_2_ net86 net97 cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1_ net367 sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_1__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput180 net180 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__343
+ VGND VGND VPWR VPWR net343 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__343/LO
+ sky130_fd_sc_hd__conb_1
Xoutput191 net191 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output281_A net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1__367 VGND VGND VPWR VPWR net367 sb_1__1_.mux_bottom_track_37.mux_l2_in_1__367/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_3__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_0__A0 sb_1__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__324__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput71 chany_bottom_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xinput82 chany_bottom_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_21.ccff_tail net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
Xinput93 chany_top_in_0[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net338 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3_ net297 net119 cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_5.mux_l1_in_2_ net83 net60 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_6.mux_l2_in_3__404 VGND VGND VPWR VPWR net404 sb_1__1_.mux_top_track_6.mux_l2_in_3__404/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_3__S sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chanx_right_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__330
+ VGND VGND VPWR VPWR net330 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__330/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_2_ net27 net8 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold29_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_15.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X net148 VGND VGND VPWR VPWR
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_59_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__319__A sb_1__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_2__A0 sb_1__1_.mux_left_track_13.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_2__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_2__A0 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l2_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input88_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l2_in_3_ net385 net26 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_48_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_10.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_2__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_1__S sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_4__A0 sb_1__1_.mux_left_track_45.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input142_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_24_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_0.mux_l4_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_2__S sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.mux_l3_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.ccff_head VGND
+ VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_1.ccff_head
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ net439 VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net340 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__mux2_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_0__S sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__332__A sb_1__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_20.mux_l1_in_1_ net36 net41 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ net76 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_289_ sb_1__1_.mux_right_track_36.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3_ net308 net104 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_64_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__327__A sb_1__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_0__A0 sb_1__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__355
+ VGND VGND VPWR VPWR net355 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__355/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_45.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l4_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_2_ net31 net39 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input105_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_1__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_53.mux_l2_in_1_ net381 sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_1__S sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_52.mux_l2_in_1__403 VGND VGND VPWR VPWR net403 sb_1__1_.mux_top_track_52.mux_l2_in_1__403/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_1_ net66 cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_10.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_2__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l2_in_3_ net397 net3 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output274_A net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_3__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_12.mux_l3_in_1_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 chany_bottom_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput94 chany_top_in_0[10] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xinput83 chany_bottom_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__340__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_5.mux_l1_in_1_ net47 net117 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.mux_l1_in_2_ net283 net87 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_37.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_5.mux_l4_in_0_ net438 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X
+ cby_1__1_.mem_right_ipin_5.ccff_tail VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__250__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input33_A chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_1__S sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_1_ net270 net38 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_5_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_39_prog_clk net469 net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_3__S sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__335__A sb_1__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_1__S sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_0__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_12.mux_l2_in_2_ net12 net86 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_11.mux_l2_in_3_ net373 net285 sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_2.mux_l4_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_10.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_1_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ net437 cby_1__1_.mem_right_ipin_5.mem_out\[2\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_4__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input135_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_5_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3__412 VGND VGND VPWR VPWR net412 cbx_1__1_.mux_top_ipin_15.mux_l2_in_3__412/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_2__A0 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_20.mux_l1_in_0_ net140 net142 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_4_ net281 net279 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_2.mux_l3_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_357_ sb_1__1_.mux_top_track_20.out VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_288_ net5 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_2_ net63 net94 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XFILLER_64_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_44.mux_l3_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net354 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__343__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_45.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_4__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l4_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA__253__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_53.mux_l2_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_1__A0 net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_4.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_10.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_2__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_3__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_1__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_1__S sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__338__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_0__A0 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_52_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_5.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput160 net160 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput193 net193 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_2.mux_l2_in_2_ net32 net18 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__248__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_2__S cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_1_ net402 sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_12.mux_l3_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3__409 VGND VGND VPWR VPWR net409 cbx_1__1_.mux_top_ipin_12.mux_l2_in_3__409/LO
+ sky130_fd_sc_hd__conb_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput73 chany_bottom_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput95 chany_top_in_0[11] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3__311 VGND VGND VPWR VPWR net311 cby_1__1_.mux_right_ipin_8.mux_l2_in_3__311/LO
+ sky130_fd_sc_hd__conb_1
Xinput84 chany_bottom_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
XFILLER_88_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net356 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l3_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_29_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_53.mux_l1_in_1_ net65 net35 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_4__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_0__A0 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l1_in_0__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_0_ net53 net98 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_32_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__351__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_1__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_44.mux_l1_in_2_ net7 net22 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_43_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__352
+ VGND VGND VPWR VPWR net352 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__352/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__261__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l2_in_1_ net72 sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3__362 VGND VGND VPWR VPWR net362 sb_1__1_.mux_bottom_track_11.mux_l2_in_3__362/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_2__A0 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_11.mux_l2_in_2_ net283 sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_10.ccff_head
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__346__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_2__A0 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input128_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_2__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__256__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input93_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3__308 VGND VGND VPWR VPWR net308 cby_1__1_.mux_right_ipin_5.mux_l2_in_3__308/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_13.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCD
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l1_in_2_ net79 net131 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_1__A0 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net322 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__mux2_2
XFILLER_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_11.mux_l1_in_3_ net88 net73 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_2.mux_l3_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
X_356_ net73 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_287_ net4 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_2__S sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_1_ net92 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_0__A0 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk net465
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_4__A1 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_0__S sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input56_A chanx_right_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_2__S sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_339_ net85 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_4.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_29_prog_clk sb_1__1_.mem_top_track_10.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_84_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_3__A0 sb_1__1_.mux_left_track_29.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_0__A0 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_0__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__354__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput161 net161 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput194 net194 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_1__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input110_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__264__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_3__380 VGND VGND VPWR VPWR net380 sb_1__1_.mux_left_track_5.mux_l2_in_3__380/LO
+ sky130_fd_sc_hd__conb_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_4.mux_l2_in_3_ net390 net30 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold64_A sc_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput63 net436 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput96 chany_top_in_0[12] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 chany_bottom_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
Xinput85 chany_bottom_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_11.mux_l3_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_53.mux_l1_in_0_ net95 net113 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3_ net405 net59 cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_87_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_2
XANTENNA__259__A sb_1__1_.mux_left_track_37.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_32_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3_ net361 net4 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3_ net364 net25 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_0__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_44.mux_l1_in_1_ net67 net33 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l2_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_2__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l2_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_54_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_2__A1 net279 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_3__S sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_2__S sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_2__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__313
+ VGND VGND VPWR VPWR net313 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__313/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l4_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_70_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input86_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__272__A sb_1__1_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1__D cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_11.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__345
+ VGND VGND VPWR VPWR net345 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__345/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_1__S sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l1_in_1_ net125 net116 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input140_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_1.mux_l4_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__267__A sb_1__1_.mux_left_track_21.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l1_in_2_ net80 net58 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_355_ net72 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_286_ net32 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l4_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_0__A0 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 net458 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XFILLER_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_0__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3_ net292 net44 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l3_in_1_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_67_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_0__A0 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3__293 VGND VGND VPWR VPWR net293 cbx_1__1_.mux_top_ipin_6.mux_l2_in_3__293/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net351 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__mux2_2
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_0__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A chanx_right_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net74 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_269_ net47 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_10.ccff_head
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_4.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_0__S sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_0__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xoutput151 net151 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xoutput162 net162 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
Xoutput173 net173 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_3__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input103_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_1_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__280__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_2__A0 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__A0 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_2_ net17 net90 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput64 net453 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
Xinput97 chany_top_in_0[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
Xinput75 chany_bottom_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput86 chany_bottom_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCD
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net335 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_4.mux_l2_in_3__401 VGND VGND VPWR VPWR net401 sb_1__1_.mux_top_track_4.mux_l2_in_3__401/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__275__A sb_1__1_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output272_A net272 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_41_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_38_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_2_ net21 net23 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_2.mux_l1_in_1_ net52 net140 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_2_ net6 net11 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__325
+ VGND VGND VPWR VPWR net325 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__325/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__353
+ VGND VGND VPWR VPWR net353 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__353/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_44.mux_l1_in_0_ net37 net137 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_0__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_2__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l2_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_77_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_4_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_0__S sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input79_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_0__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_3_ net273 net270 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_3_ net372 net284 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_3__S sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_12.mux_l1_in_0_ net102 net109 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_2__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0__A0
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_1_ net43 net118 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_354_ net71 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__283__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_285_ sb_1__1_.mux_right_track_44.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_0__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 net459 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_4
XFILLER_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_2_ net3 net34 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_36.mux_l3_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_4.mux_l3_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_1__S sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_2__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__278__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_1__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_268_ net46 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_2__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_2.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_2__S sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l4_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput152 net152 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_3__399 VGND VGND VPWR VPWR net399 sb_1__1_.mux_top_track_28.mux_l2_in_3__399/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_2__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input61_A chanx_right_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_3__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__348
+ VGND VGND VPWR VPWR net348 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__348/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_36.mux_l2_in_1_ net389 sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_28_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_1_ net66 sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__337
+ VGND VGND VPWR VPWR net337 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__337/LO
+ sky130_fd_sc_hd__conb_1
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xinput98 chany_top_in_0[14] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xinput65 chany_bottom_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
Xinput76 chany_bottom_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xinput87 net448 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_60_prog_clk net420
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_38_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__291__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_38_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l3_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_34_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_2.mux_l1_in_0_ net137 net142 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_1_ net274 sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_2__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__sdfrtp_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_3__A1 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_36.mux_l1_in_2_ net8 net68 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l1_in_2_ net77 net130 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__286__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk cby_1__1_.mem_right_ipin_10.ccff_head
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_2__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_2_ net275 net57 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_79_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_1.mux_l2_in_2_ net281 net278 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_95_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_2__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_2_ net276 net55 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__334
+ VGND VGND VPWR VPWR net334 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__334/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_2__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__360
+ VGND VGND VPWR VPWR net360 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__360/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net435 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_37.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input126_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l1_in_0_ net96 net103 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_353_ sb_1__1_.mux_top_track_28.out VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input91_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_284_ net30 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_1__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_1_ net32 cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_2.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_3_ net63 net64 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_2__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__349
+ VGND VGND VPWR VPWR net349 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__349/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_44.mux_l2_in_1__391 VGND VGND VPWR VPWR net391 sb_1__1_.mux_right_track_44.mux_l2_in_1__391/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__294__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ sb_1__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_267_ sb_1__1_.mux_left_track_21.out VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net324 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net333 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__mux2_4
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_2__A1 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput164 net164 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_1__S sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input54_A chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_36.mux_l2_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_42_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ sb_1__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_2__A0 sb_1__1_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput77 chany_bottom_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xinput88 chany_bottom_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xinput66 net461 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
Xinput99 chany_top_in_0[15] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_12.ccff_tail
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_3__A1 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3__304 VGND VGND VPWR VPWR net304 cby_1__1_.mux_right_ipin_15.mux_l2_in_3__304/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3_ net301 net119 cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l3_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold62_A ccff_head_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_0__S sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_36.mux_l1_in_1_ net83 net128 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_4.mux_l1_in_1_ net127 net120 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_21.mux_l2_in_3__375 VGND VGND VPWR VPWR net375 sb_1__1_.mux_left_track_21.mux_l2_in_3__375/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_1__A0 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_1__A0 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3_ net408 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_70_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_1_ net34 net51 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net319 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_2__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_1_ net41 net50 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_0__S sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_2__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3__410 VGND VGND VPWR VPWR net410 cbx_1__1_.mux_top_ipin_13.mux_l2_in_3__410/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_12.mux_l4_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_49_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_37.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_4__S sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input119_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_3__A0 net274 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ net69 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_283_ net29 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input84_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_3__A0 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_1__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_0__S sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_18_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_0__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_2_ net81 net34 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_335_ sb_1__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ net43 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__327
+ VGND VGND VPWR VPWR net327 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__327/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_3__S sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput165 net165 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_20.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A chanx_right_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk cbx_1__1_.ccff_head
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_0__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ net451 VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_318_ net95 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
X_249_ net55 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput67 chany_bottom_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
Xinput89 chany_bottom_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_4
Xinput78 chany_bottom_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3__407 VGND VGND VPWR VPWR net407 cbx_1__1_.mux_top_ipin_10.mux_l2_in_3__407/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_84_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_2__S sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input101_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_2__A0 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk sb_1__1_.mem_right_track_52.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_8.ccff_tail
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_1__S sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_3__S sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_1__A0 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_1__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_36.mux_l1_in_0_ net96 net98 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l1_in_0_ net107 net113 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_1__S sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_1__S sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output270_A net270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_3__S sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l2_in_1__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net416 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3_ net298 net118 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_50_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_3__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_2.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_1__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_2_ net26 net37 cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_1__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_0_ net94 net111 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_1__S sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_3__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_0_ net115 net101 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3__306 VGND VGND VPWR VPWR net306 cby_1__1_.mux_right_ipin_3.mux_l2_in_3__306/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold18_A test_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.ccff_tail
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_351_ net68 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_3__A1 net271 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_282_ net28 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_45.mux_l3_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_1__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_3__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output233_A net233 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.ccff_tail
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_1.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_1.mux_l1_in_1_ net51 net94 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_2__A0 sb_1__1_.mux_left_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input131_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l4_in_0_ net450 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ cby_1__1_.mem_right_ipin_1.ccff_tail VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_334_ sb_1__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ net42 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_3__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l2_in_2__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput166 net166 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
XFILLER_95_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1_ net368 sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_20.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_1__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net315 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__mux2_2
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_317_ net94 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3_ net309 net119 cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
X_248_ net44 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput68 chany_bottom_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput79 chany_bottom_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_0__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_0__S sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_1__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net360 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net147 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_1_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ net449 cby_1__1_.mem_right_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_52.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_0__S sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_40_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_2_ net3 net7 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_hold48_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l1_in_0__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_1__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_1__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_88_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_37_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 net418 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_right_track_20.mux_l2_in_3_ net387 net25 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_94_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_2_ net87 net98 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_5.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ net446 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_2.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l4_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_1__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_1_ net6 cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net337 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_3__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_0__S sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_52.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ net67 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_281_ sb_1__1_.mux_right_track_52.out VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_3__S sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_1.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_1.mux_l1_in_0_ net111 net114 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_2__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3__291 VGND VGND VPWR VPWR net291 cbx_1__1_.mux_top_ipin_4.mux_l2_in_3__291/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_20.mux_l4_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_58_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_3__S sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_333_ net111 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_264_ net41 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_0__A0 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__316
+ VGND VGND VPWR VPWR net316 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__316/LO
+ sky130_fd_sc_hd__conb_1
Xoutput167 net167 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput156 net156 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
XFILLER_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_20.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_316_ net122 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_4
Xinput14 net442 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput69 chany_bottom_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_0__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_20.mux_l3_in_1_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_8.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_2__A0 net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_87_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_44.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_7.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_27_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_A chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_78_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ net452 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_40_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_3__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_1_ net271 net37 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_3__396 VGND VGND VPWR VPWR net396 sb_1__1_.mux_top_track_12.mux_l2_in_3__396/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_1.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__319
+ VGND VGND VPWR VPWR net319 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__319/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_20.mux_l2_in_2_ net11 net85 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xhold3 prog_reset VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_1_ net67 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold60_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_2.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_0__S sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_20.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_21.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_1__S sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_60_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_52.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_280_ net26 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk net472 net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_1__S sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_1__A0 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l2_in_3_ net383 net4 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_1.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold23_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_52.mux_l3_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_0__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_2__S sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_3__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input117_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ sb_1__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_0__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_263_ sb_1__1_.mux_left_track_29.out VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input82_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput168 net168 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
XANTENNA__303__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 net179 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_0__A0 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_12.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_45.mux_l2_in_1__379 VGND VGND VPWR VPWR net379 sb_1__1_.mux_left_track_45.mux_l2_in_1__379/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_315_ sb_1__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_56_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_4
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_52.mux_l2_in_1_ net403 sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_20.mux_l3_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_2__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_3__S sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_7.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l4_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A chanx_right_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_0_ net54 net97 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_0__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_52.mux_l1_in_2_ net5 net23 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_2__S sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_1_ net71 sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__335
+ VGND VGND VPWR VPWR net335 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__335/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 net414 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_2__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3_ net406 net58 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_0.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__311__A sb_1__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_3__S sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk sb_1__1_.mem_top_track_20.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_65_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l3_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_70_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_2__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_1__S sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net341 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net355 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_29.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_2__S sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_10.mux_l2_in_3_ net395 net28 sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_44.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_53.mux_l1_in_0__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.mux_l1_in_2_ net80 net132 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_29.mux_l2_in_3_ net376 net280 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_76_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net326 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_2_ net21 net87 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__1_.mem_bottom_track_53.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_1__S cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_3__A1 net284 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_331_ sb_1__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_262_ net39 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_input75_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_1__S sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l1_in_4_ net13 net88 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput158 net158 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
XFILLER_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_2_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_31_prog_clk cby_1__1_.ccff_tail net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_2__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_314_ net120 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_2__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output279_A net279 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_52.mux_l2_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_10.mux_l4_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3_ net293 net59 cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_2__A0 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.mux_l4_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA__314__A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net352 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__mux2_2
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_7.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3_ net371 net29 sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3__302 VGND VGND VPWR VPWR net302 cby_1__1_.mux_right_ipin_13.mux_l2_in_3__302/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input38_A chanx_right_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_2__S sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__309__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_1__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_10.mux_l3_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_52.mux_l1_in_1_ net65 net35 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_6.mux_l2_in_3__393 VGND VGND VPWR VPWR net393 sb_1__1_.mux_right_track_6.mux_l2_in_3__393/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_94_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 net123 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_2__S sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l3_in_1_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_61_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_2__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold46_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_4__S cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_2_ net27 net38 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_12.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l3_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_65_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_4_ net19 net273 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_3__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_1__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_3__A1 net285 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_2__S sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_7.mux_l4_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_2_ net6 sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__322__A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[2\] net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_36_prog_clk_A clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_20.mux_l1_in_1_ net126 net115 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l2_in_2_ net74 net69 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_1__S sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3__297 VGND VGND VPWR VPWR net297 cby_1__1_.mux_right_ipin_0.mux_l2_in_3__297/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__342
+ VGND VGND VPWR VPWR net342 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__342/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l2_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_82_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__317__A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_2__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ net108 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ net38 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_0__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input68_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_12.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_2__S sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_10.mux_l1_in_3_ net73 net58 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput148 net148 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XFILLER_87_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_1__S sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_2__A0 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input122_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l1_in_2_ net131 net128 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_42_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_313_ net119 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_8
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_2__S sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_44.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_2__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_0__S sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3__406 VGND VGND VPWR VPWR net406 cbx_1__1_.mux_top_ipin_1.mux_l2_in_3__406/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_1__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__330__A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_5.ccff_tail
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_3__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_2_ net16 sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net330 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_4__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_60_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__325__A net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l3_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_52.mux_l1_in_0_ net54 net138 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input50_A chanx_right_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 net473 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_29.mux_l3_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_61_prog_clk net463 net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_2__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l2_in_2__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_1_ net7 cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_26_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_3_ net271 net269 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_3_ net382 net284 sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_4.mux_l1_in_3__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_21.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input98_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_load_slew288_A net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_20.mux_l1_in_0_ net101 net105 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_30_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__321
+ VGND VGND VPWR VPWR net321 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__321/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_2__S sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_29.mux_l2_in_1_ net70 net44 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_0.mux_l2_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net344 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_4_ net280 net278 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_82_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3__371 VGND VGND VPWR VPWR net371 sb_1__1_.mux_bottom_track_7.mux_l2_in_3__371/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_6.mux_l2_in_1__S sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__333__A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_44.mux_l3_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_3__A0 net272 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_20.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_260_ net37 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_12.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_7.mux_l4_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_60_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l1_in_2_ net43 net45 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput149 net149 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__1_.mux_right_ipin_1.mux_l2_in_2__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_1__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_29_prog_clk sb_1__1_.mem_right_track_0.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__328__A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk sb_1__1_.mem_bottom_track_1.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_74_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_0__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input115_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l1_in_1_ net125 net93 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_312_ net118 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input80_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_44.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_bottom_track_45.mux_l1_in_2__S sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_44.mux_l2_in_1_ net391 sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l2_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_1__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_87_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_20.mux_l2_in_3__387 VGND VGND VPWR VPWR net387 sb_1__1_.mux_right_track_20.mux_l2_in_3__387/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mux_right_ipin_12.mux_l1_in_3__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l1_in_0__A1 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_2__A0 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output284_A net284 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net334 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__mux2_4
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_55_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_12.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__251__A sb_1__1_.mux_left_track_53.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_44.mux_l1_in_2_ net7 net67 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A chanx_right_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 net1 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_2__S sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_2_ net275 net59 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_7.mux_l2_in_2_ net282 sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__336__A sb_1__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_12.mux_l2_in_2__S sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_1__A0 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3_ net302 net115 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_44.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_0__S cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l1_in_1__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[0\] net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.mux_l2_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_3__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_7.mux_l1_in_3_ net89 net76 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3_ net409 net59 cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_3__A1 net270 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_12.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_10.mux_l1_in_1_ net140 net138 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_13.mux_l4_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_0.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.mux_l1_in_1_ net39 net104 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__344__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_1__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input108_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_0.mux_l1_in_0_ net94 net111 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
X_311_ sb_1__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_4
XANTENNA__254__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_36.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_input73_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_44.mux_l2_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_2__S sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_2__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_2__S sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__339__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_4__A0 sb_1__1_.mux_left_track_37.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__249__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_3.mux_l1_in_2__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l2_in_3__S cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_1_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_0__S sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_1__S sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3__296 VGND VGND VPWR VPWR net296 cbx_1__1_.mux_top_ipin_9.mux_l2_in_3__296/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_1_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_12.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_6.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_44.mux_l1_in_1_ net84 net129 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 net475 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input36_A chanx_right_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_0__S sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l2_in_3__A1 sb_1__1_.mux_left_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l2_in_1__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l1_in_1__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_0__A0 sb_1__1_.mux_left_track_3.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_1_ net40 net46 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__352__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_2
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_4.mux_l1_in_1__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_2_ net74 net95 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_44_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_44.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__262__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_head net289 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__347__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_4__S sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input138_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_3__A1 net284 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA__257__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_3_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l1_in_3__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3_ net305 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_2_ net82 net59 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_4__A0 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_10.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_10.mux_l1_in_0_ net136 net142 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_3__S sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l2_in_1__A0 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk net464 net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_right_track_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__1_.mux_top_ipin_8.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_29.mux_l1_in_0_ net99 net109 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_7__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__360__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_2__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_2.mux_l2_in_1__S sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_0__S sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_310_ net116 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_1__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__270__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0__A1
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_3.mux_l2_in_3__S sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_1__402 VGND VGND VPWR VPWR net402 sb_1__1_.mux_top_track_44.mux_l2_in_1__402/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_5.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__355__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l4_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_78_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input120_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__265__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_0_ net454 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mem_right_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_10.mux_l2_in_3__395 VGND VGND VPWR VPWR net395 sb_1__1_.mux_top_track_10.mux_l2_in_3__395/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ net457 VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_1__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l2_in_3__376 VGND VGND VPWR VPWR net376 sb_1__1_.mux_left_track_29.mux_l2_in_3__376/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_4.mux_l2_in_3__390 VGND VGND VPWR VPWR net390 sb_1__1_.mux_right_track_4.mux_l2_in_3__390/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_top_track_12.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_6.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net316 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__mux2_4
Xsb_1__1_.mux_right_track_44.mux_l1_in_0_ net121 net97 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3_ net310 sb_1__1_.mux_bottom_track_45.out cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xhold9 net2 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_1_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_11_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_6.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_0_ net119 net106 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_0__A0 sb_1__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_1__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_1_ net64 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_36.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_38_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR cby_1__1_.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_1__1_.mux_right_ipin_3.mux_l2_in_3__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l2_in_3_ net401 net27 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_11.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__363__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_1__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_top_track_20.mux_l2_in_3__S sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input96_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__273__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_53.mux_l3_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_53.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_25_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_7.mux_l1_in_1_ net46 net119 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_load_slew286_A net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_7.mux_l4_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l1_in_4__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_2_ net101 net70 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__358__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_2__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_2__S sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_1__A1 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__268__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_right_track_0.ccff_head
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l2_in_1__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1_ net370 sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_2__A0 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_13.mux_l2_in_3_ net374 net284 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_4.mux_l4_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_1__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mux_right_ipin_14.mux_l2_in_3__A1 sb_1__1_.mux_bottom_track_53.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_1_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_60_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_1__S sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_2__A0 net280 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__A0 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3__300 VGND VGND VPWR VPWR net300 cby_1__1_.mux_right_ipin_11.mux_l2_in_3__300/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input113_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_2_ net5 net24 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_28.mux_l2_in_1__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l3_in_1_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_17_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__1_.mux_top_track_4.mux_l2_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_2__A0 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_30_prog_clk sb_1__1_.mem_right_track_6.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_29_prog_clk sb_1__1_.mem_top_track_10.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xoutput280 net280 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_2_ net90 net101 cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_59_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__276__A sb_1__1_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_output282_A net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_53_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_0__S sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l4_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__317
+ VGND VGND VPWR VPWR net317 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__317/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_88_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net345 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__mux2_4
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_37_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_15_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input41_A chanx_right_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_1__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3_ net362 net28 sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_54_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_4.mux_l2_in_2_ net30 net17 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l2_in_1__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_2__A0 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_1__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l1_in_1__S sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input89_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_0_ net121 net106 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l3_in_1_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_13.mux_l2_in_3__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net432 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_2__A0 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_right_track_36.mux_l1_in_2__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_4_ net15 net274 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net347 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__284__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_36.mem_out\[1\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_11.mux_l4_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_86_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_11.mux_l2_in_2__S sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_13.mux_l2_in_2_ net278 net86 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_37.mux_l1_in_2__A1 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__357
+ VGND VGND VPWR VPWR net357 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__357/LO
+ sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ net455 VGND VGND VPWR VPWR
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_2__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__279__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_33_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_368_ net146 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_299_ net17 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_1__A0 sb_1__1_.mux_left_track_7.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold12_A reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l2_in_3__S sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l1_in_0__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_2__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_6.mux_l1_in_2__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_1.mux_l2_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_1_1__f_clk0_A clknet_0_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input106_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input71_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_0__A0 sb_1__1_.mux_left_track_1.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__S sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_61_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_1_ net272 net33 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l3_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_11.mux_l1_in_2__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_4.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_1_ net70 cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput270 net270 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
Xoutput281 net281 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
XFILLER_58_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_0__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__292__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output275_A net275 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_0__A0 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_0__A0 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_21.mux_l2_in_3__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A chanx_right_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_1.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3__312 VGND VGND VPWR VPWR net312 cby_1__1_.mux_right_ipin_9.mux_l2_in_3__312/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_2_ net13 sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__287__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_0_prog_clk_A clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_4.mux_l2_in_1_ net90 sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_2__A0 net283 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_right_track_44.mux_l1_in_2__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_61_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_4.mux_l2_in_3__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_head
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_2__A0 net276 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_3_ net393 net29 sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_0__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_2__A0 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_28.mux_l1_in_0__A1 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l3_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3_ net413 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_45.mux_l1_in_2__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_47_prog_clk cby_1__1_.mem_right_ipin_11.ccff_tail
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__324
+ VGND VGND VPWR VPWR net324 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__324/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_3_ net272 net270 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input136_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3_ net366 net32 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_66_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_4.mux_l1_in_2_ net77 net60 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_36.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_4_ net89 net70 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_35_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3__377 VGND VGND VPWR VPWR net377 sb_1__1_.mux_left_track_3.mux_l2_in_3__377/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ net460 VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_13.mux_l2_in_1_ net72 sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_7.mux_l2_in_2__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_3__S sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3__309 VGND VGND VPWR VPWR net309 cby_1__1_.mux_right_ipin_6.mux_l2_in_3__309/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__295__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3__364 VGND VGND VPWR VPWR net364 sb_1__1_.mux_bottom_track_21.mux_l2_in_3__364/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_367_ sb_1__1_.mux_top_track_0.out VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ net16 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_6.mux_l4_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_2__S sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_34_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk net462
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_0_ net35 net95 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l4_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_13.mux_l1_in_2_ net79 net56 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_0__A0 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xoutput260 net260 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput271 net271 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xoutput282 net282 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
XFILLER_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3_ net294 sb_1__1_.mux_left_track_45.out cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_70_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_12.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_right_track_52.mux_l1_in_2__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l3_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_36.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_1__S sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_0__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_3__A0 sb_1__1_.mux_bottom_track_29.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_4__A0 net280 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_46_prog_clk cby_1__1_.mem_right_ipin_14.ccff_tail
+ net415 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__1_.mux_top_track_36.mux_l1_in_0__A1 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_90_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_13.mux_l2_in_2__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l2_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net336 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_53.mux_l1_in_2__A1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net327 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__mux2_4
XFILLER_93_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_2__A0 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_0__S sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__RESET_B
+ net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_3.mux_l1_in_2__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_2_ net16 sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l1_in_4__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l1_in_0__A1 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_10.mux_l1_in_2__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__298__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net432 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_2.mux_l1_in_1__S sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l2_in_2__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_1__A0 sb_1__1_.mux_bottom_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold35_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_7.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_2_ net276 net58 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_2_ net18 net22 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XANTENNA_input129_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_72_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_4.mux_l1_in_1_ net47 net50 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4__f_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input94_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_sb_1__1_.mux_left_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_1__S sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_28.ccff_tail
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_63_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_7.ccff_tail
+ net286 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_0_clk0_A clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_1__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_48_prog_clk net468 net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_3_ net76 net131 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_24_prog_clk_A clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_13.mux_l2_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__346
+ VGND VGND VPWR VPWR net346 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__346/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_366_ sb_1__1_.mux_top_track_2.out VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ sb_1__1_.mux_right_track_20.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__1_.mux_top_track_52.mux_l1_in_0__A0 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_7.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_3_ net274 net271 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3_ net377 net285 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_11.mux_l1_in_4__S sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l2_in_3__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net325 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[2\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input57_A chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_2__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_349_ sb_1__1_.mux_top_track_36.out VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3__294 VGND VGND VPWR VPWR net294 cbx_1__1_.mux_top_ipin_7.mux_l2_in_3__294/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l1_in_1_ net42 net116 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mux_top_track_44.mux_l1_in_0__A1 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput250 net250 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput261 net261 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput283 net283 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput272 net272 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input111_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_2_ net30 net41 cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] net287 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l3_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_36.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_29.mux_l2_in_2__S sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_top_track_10.mux_l1_in_0__A0 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_1.ccff_tail
+ net288 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_2.mux_l1_in_3__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_4__A1 net278 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_right_track_0.mux_l1_in_2__S sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_90_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_6.mux_l2_in_2__S sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l4_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XANTENNA_output280_A net280 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_5.mux_l2_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_1__1_.mux_right_ipin_0.mux_l1_in_4__S cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_6.mux_l2_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_80_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_5.mux_l2_in_2__S sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold60 ccff_head_1 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_1__1_.mux_right_ipin_15.mux_l1_in_1__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_7.mux_l2_in_3__A1 net284 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_14_prog_clk_A clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_1_ net43 net45 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_53_prog_clk_A clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l3_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_2__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_82_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l1_in_0_ net138 net135 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_1__A0 sb_1__1_.mux_left_track_11.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_3_ net399 net14 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_56_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_2_ net129 net127 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_3__372 VGND VGND VPWR VPWR net372 sb_1__1_.mux_left_track_1.mux_l2_in_3__372/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input141_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_365_ sb_1__1_.mux_top_track_4.out VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_296_ net13 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_2_ net276 net61 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_1__A0 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_3.mux_l2_in_2_ net282 net279 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_4.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_55_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_52_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[2\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_348_ net65 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_1__1_.mux_right_ipin_13.mux_l2_in_2__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_279_ net25 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_1.mux_l1_in_1__S sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_13.mux_l1_in_0_ net100 net102 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0__CLK
+ clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__350
+ VGND VGND VPWR VPWR net350 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__350/LO
+ sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__339
+ VGND VGND VPWR VPWR net339 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__339/LO
+ sky130_fd_sc_hd__conb_1
Xoutput240 net240 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput251 net251 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput262 net262 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_28.mux_l4_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xoutput284 net284 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
XFILLER_58_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput273 net273 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_1_ net10 cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input104_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_34_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[0\] net287 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mux_top_track_10.mux_l2_in_1__S sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__1_.mem_top_track_28.ccff_tail
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_37.mux_l3_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_3.mux_l1_in_3_ net92 net78 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_1__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0__SCE
+ net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output273_A net273 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_13.mux_l2_in_3__374 VGND VGND VPWR VPWR net374 sb_1__1_.mux_left_track_13.mux_l2_in_3__374/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_2__A0 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_28.mux_l3_in_1_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_2__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_43_prog_clk_A clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_25_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net287 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_6.mux_l2_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_9.mux_l2_in_3__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_37.mux_l2_in_1_ net378 sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_41_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold50 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold61 net419 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_0__A0 sb_1__1_.mux_bottom_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_0__A0 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l3_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_0_ net118 net103 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_28.mem_out\[2\]
+ net289 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3_ net303 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_left_track_21.mux_l1_in_1__S sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net415 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_2__A0 net278 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l3_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_17_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_7.ccff_tail
+ net286 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_top_track_28.mux_l2_in_2__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__1_.mux_top_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_4.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_28.mux_l2_in_2_ net9 net19 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xinput140 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_2__A0 sb_1__1_.mux_bottom_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold40_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l1_in_1_ net125 net119 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net317 net430 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_37.mux_l1_in_2_ net281 net66 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_26_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_364_ sb_1__1_.mux_top_track_6.out VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
X_295_ net12 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l2_in_1__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XANTENNA_cbx_1__1_.mux_top_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_52.mux_l2_in_1_ net392 sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3_ net410 net55 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_51_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_bottom_track_7.mux_l1_in_1__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_1_ net62 net48 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_1__1_.mux_right_ipin_4.mux_l1_in_4__A0 sb_1__1_.mux_bottom_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net343 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_39_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net289 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[0\] net288 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[1\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_15.mux_l2_in_3__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
X_347_ net64 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_278_ net14 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_14.mux_l4_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__1_.mux_top_ipin_14.mux_l1_in_0__A0 sb_1__1_.mux_left_track_5.out VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3__299 VGND VGND VPWR VPWR net299 cby_1__1_.mux_right_ipin_10.mux_l2_in_3__299/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_83_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net415 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput241 net241 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput252 net252 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput230 net230 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput285 net285 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput263 net263 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput274 net274 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_left_track_7.mux_l1_in_0__S sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk
+ sb_1__1_.mem_bottom_track_45.ccff_tail net287 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net314 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chanx_right_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_52.mux_l1_in_2_ net5 net63 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8__RESET_B
+ net289 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_2_ net84 net62 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_bottom_track_29.mux_l2_in_1__A0 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_20.mux_l2_in_2__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net287 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_prog_clk_A clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_12.mux_l1_in_2__A0 sb_1__1_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_1__1_.mux_right_ipin_10.mux_l1_in_1__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l4_in_0_ net444 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X
+ cbx_1__1_.mem_top_ipin_13.ccff_tail VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__D sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__1_.mux_left_track_1.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net288 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__1_.mux_bottom_track_5.mux_l2_in_2__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_28.mux_l3_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_91_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_left_track_21.mux_l2_in_2__A0 net279 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_right_track_12.mux_l2_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_1__S sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l2_in_3_ net384 net28 sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__1_.mux_top_ipin_10.mux_l1_in_4__A0 sb_1__1_.mux_left_track_45.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__D sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_37.mux_l2_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 chany_bottom_in[10] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold62 ccff_head_2 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold51 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1__368 VGND VGND VPWR VPWR net368 sb_1__1_.mux_bottom_track_45.mux_l2_in_1__368/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mux_right_ipin_8.mux_l1_in_0__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_4 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_cbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net288 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__1_.mux_top_track_0.mux_l1_in_0__A1 net141 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_53.mux_l2_in_1__381 VGND VGND VPWR VPWR net381 sb_1__1_.mux_left_track_53.mux_l2_in_1__381/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__1_.mux_top_track_2.mux_l2_in_2__S sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__1_.mux_top_ipin_9.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk net471 net286 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net289 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14__RESET_B
+ net415 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_28.mem_out\[1\]
+ net288 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ net443 cbx_1__1_.mem_top_ipin_13.mem_out\[2\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__1_.mux_left_track_13.mux_l2_in_2__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__1_.mux_right_track_0.mux_l2_in_0__S sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.mem_out\[0\]
+ net287 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l2_in_1_ net74 net69 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput130 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xinput141 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net141 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__1_.mux_left_track_1.mux_l2_in_2__S sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net288 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__347
+ VGND VGND VPWR VPWR net347 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__347/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cby_1__1_.mux_right_ipin_6.mux_l1_in_2__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mux_bottom_track_37.mux_l1_in_2__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net287 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_10.mux_l1_in_4_ net88 net73 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_right_track_6.mux_l1_in_0_ net106 net112 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net286 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

