magic
tech sky130A
magscale 1 2
timestamp 1656943670
<< viali >>
rect 2881 4573 2915 4607
rect 9229 4573 9263 4607
rect 2513 3893 2547 3927
rect 3709 3893 3743 3927
rect 7757 3893 7791 3927
rect 9045 3893 9079 3927
rect 2697 3485 2731 3519
rect 9229 3485 9263 3519
<< metal1 >>
rect 1104 11450 10856 11472
rect 1104 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 2302 11450
rect 2354 11398 2366 11450
rect 2418 11398 2430 11450
rect 2482 11398 4622 11450
rect 4674 11398 4686 11450
rect 4738 11398 4750 11450
rect 4802 11398 4814 11450
rect 4866 11398 4878 11450
rect 4930 11398 7070 11450
rect 7122 11398 7134 11450
rect 7186 11398 7198 11450
rect 7250 11398 7262 11450
rect 7314 11398 7326 11450
rect 7378 11398 9518 11450
rect 9570 11398 9582 11450
rect 9634 11398 9646 11450
rect 9698 11398 9710 11450
rect 9762 11398 9774 11450
rect 9826 11398 10856 11450
rect 1104 11376 10856 11398
rect 1104 10906 10856 10928
rect 1104 10854 3398 10906
rect 3450 10854 3462 10906
rect 3514 10854 3526 10906
rect 3578 10854 3590 10906
rect 3642 10854 3654 10906
rect 3706 10854 5846 10906
rect 5898 10854 5910 10906
rect 5962 10854 5974 10906
rect 6026 10854 6038 10906
rect 6090 10854 6102 10906
rect 6154 10854 8294 10906
rect 8346 10854 8358 10906
rect 8410 10854 8422 10906
rect 8474 10854 8486 10906
rect 8538 10854 8550 10906
rect 8602 10854 10856 10906
rect 1104 10832 10856 10854
rect 1104 10362 10856 10384
rect 1104 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 2302 10362
rect 2354 10310 2366 10362
rect 2418 10310 2430 10362
rect 2482 10310 4622 10362
rect 4674 10310 4686 10362
rect 4738 10310 4750 10362
rect 4802 10310 4814 10362
rect 4866 10310 4878 10362
rect 4930 10310 7070 10362
rect 7122 10310 7134 10362
rect 7186 10310 7198 10362
rect 7250 10310 7262 10362
rect 7314 10310 7326 10362
rect 7378 10310 9518 10362
rect 9570 10310 9582 10362
rect 9634 10310 9646 10362
rect 9698 10310 9710 10362
rect 9762 10310 9774 10362
rect 9826 10310 10856 10362
rect 1104 10288 10856 10310
rect 1104 9818 10856 9840
rect 1104 9766 3398 9818
rect 3450 9766 3462 9818
rect 3514 9766 3526 9818
rect 3578 9766 3590 9818
rect 3642 9766 3654 9818
rect 3706 9766 5846 9818
rect 5898 9766 5910 9818
rect 5962 9766 5974 9818
rect 6026 9766 6038 9818
rect 6090 9766 6102 9818
rect 6154 9766 8294 9818
rect 8346 9766 8358 9818
rect 8410 9766 8422 9818
rect 8474 9766 8486 9818
rect 8538 9766 8550 9818
rect 8602 9766 10856 9818
rect 1104 9744 10856 9766
rect 1104 9274 10856 9296
rect 1104 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 2302 9274
rect 2354 9222 2366 9274
rect 2418 9222 2430 9274
rect 2482 9222 4622 9274
rect 4674 9222 4686 9274
rect 4738 9222 4750 9274
rect 4802 9222 4814 9274
rect 4866 9222 4878 9274
rect 4930 9222 7070 9274
rect 7122 9222 7134 9274
rect 7186 9222 7198 9274
rect 7250 9222 7262 9274
rect 7314 9222 7326 9274
rect 7378 9222 9518 9274
rect 9570 9222 9582 9274
rect 9634 9222 9646 9274
rect 9698 9222 9710 9274
rect 9762 9222 9774 9274
rect 9826 9222 10856 9274
rect 1104 9200 10856 9222
rect 1104 8730 10856 8752
rect 1104 8678 3398 8730
rect 3450 8678 3462 8730
rect 3514 8678 3526 8730
rect 3578 8678 3590 8730
rect 3642 8678 3654 8730
rect 3706 8678 5846 8730
rect 5898 8678 5910 8730
rect 5962 8678 5974 8730
rect 6026 8678 6038 8730
rect 6090 8678 6102 8730
rect 6154 8678 8294 8730
rect 8346 8678 8358 8730
rect 8410 8678 8422 8730
rect 8474 8678 8486 8730
rect 8538 8678 8550 8730
rect 8602 8678 10856 8730
rect 1104 8656 10856 8678
rect 1104 8186 10856 8208
rect 1104 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 2302 8186
rect 2354 8134 2366 8186
rect 2418 8134 2430 8186
rect 2482 8134 4622 8186
rect 4674 8134 4686 8186
rect 4738 8134 4750 8186
rect 4802 8134 4814 8186
rect 4866 8134 4878 8186
rect 4930 8134 7070 8186
rect 7122 8134 7134 8186
rect 7186 8134 7198 8186
rect 7250 8134 7262 8186
rect 7314 8134 7326 8186
rect 7378 8134 9518 8186
rect 9570 8134 9582 8186
rect 9634 8134 9646 8186
rect 9698 8134 9710 8186
rect 9762 8134 9774 8186
rect 9826 8134 10856 8186
rect 1104 8112 10856 8134
rect 1104 7642 10856 7664
rect 1104 7590 3398 7642
rect 3450 7590 3462 7642
rect 3514 7590 3526 7642
rect 3578 7590 3590 7642
rect 3642 7590 3654 7642
rect 3706 7590 5846 7642
rect 5898 7590 5910 7642
rect 5962 7590 5974 7642
rect 6026 7590 6038 7642
rect 6090 7590 6102 7642
rect 6154 7590 8294 7642
rect 8346 7590 8358 7642
rect 8410 7590 8422 7642
rect 8474 7590 8486 7642
rect 8538 7590 8550 7642
rect 8602 7590 10856 7642
rect 1104 7568 10856 7590
rect 1104 7098 10856 7120
rect 1104 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 2302 7098
rect 2354 7046 2366 7098
rect 2418 7046 2430 7098
rect 2482 7046 4622 7098
rect 4674 7046 4686 7098
rect 4738 7046 4750 7098
rect 4802 7046 4814 7098
rect 4866 7046 4878 7098
rect 4930 7046 7070 7098
rect 7122 7046 7134 7098
rect 7186 7046 7198 7098
rect 7250 7046 7262 7098
rect 7314 7046 7326 7098
rect 7378 7046 9518 7098
rect 9570 7046 9582 7098
rect 9634 7046 9646 7098
rect 9698 7046 9710 7098
rect 9762 7046 9774 7098
rect 9826 7046 10856 7098
rect 1104 7024 10856 7046
rect 1104 6554 10856 6576
rect 1104 6502 3398 6554
rect 3450 6502 3462 6554
rect 3514 6502 3526 6554
rect 3578 6502 3590 6554
rect 3642 6502 3654 6554
rect 3706 6502 5846 6554
rect 5898 6502 5910 6554
rect 5962 6502 5974 6554
rect 6026 6502 6038 6554
rect 6090 6502 6102 6554
rect 6154 6502 8294 6554
rect 8346 6502 8358 6554
rect 8410 6502 8422 6554
rect 8474 6502 8486 6554
rect 8538 6502 8550 6554
rect 8602 6502 10856 6554
rect 1104 6480 10856 6502
rect 1104 6010 10856 6032
rect 1104 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 2302 6010
rect 2354 5958 2366 6010
rect 2418 5958 2430 6010
rect 2482 5958 4622 6010
rect 4674 5958 4686 6010
rect 4738 5958 4750 6010
rect 4802 5958 4814 6010
rect 4866 5958 4878 6010
rect 4930 5958 7070 6010
rect 7122 5958 7134 6010
rect 7186 5958 7198 6010
rect 7250 5958 7262 6010
rect 7314 5958 7326 6010
rect 7378 5958 9518 6010
rect 9570 5958 9582 6010
rect 9634 5958 9646 6010
rect 9698 5958 9710 6010
rect 9762 5958 9774 6010
rect 9826 5958 10856 6010
rect 1104 5936 10856 5958
rect 1104 5466 10856 5488
rect 1104 5414 3398 5466
rect 3450 5414 3462 5466
rect 3514 5414 3526 5466
rect 3578 5414 3590 5466
rect 3642 5414 3654 5466
rect 3706 5414 5846 5466
rect 5898 5414 5910 5466
rect 5962 5414 5974 5466
rect 6026 5414 6038 5466
rect 6090 5414 6102 5466
rect 6154 5414 8294 5466
rect 8346 5414 8358 5466
rect 8410 5414 8422 5466
rect 8474 5414 8486 5466
rect 8538 5414 8550 5466
rect 8602 5414 10856 5466
rect 1104 5392 10856 5414
rect 1104 4922 10856 4944
rect 1104 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 2302 4922
rect 2354 4870 2366 4922
rect 2418 4870 2430 4922
rect 2482 4870 4622 4922
rect 4674 4870 4686 4922
rect 4738 4870 4750 4922
rect 4802 4870 4814 4922
rect 4866 4870 4878 4922
rect 4930 4870 7070 4922
rect 7122 4870 7134 4922
rect 7186 4870 7198 4922
rect 7250 4870 7262 4922
rect 7314 4870 7326 4922
rect 7378 4870 9518 4922
rect 9570 4870 9582 4922
rect 9634 4870 9646 4922
rect 9698 4870 9710 4922
rect 9762 4870 9774 4922
rect 9826 4870 10856 4922
rect 1104 4848 10856 4870
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3786 4604 3792 4616
rect 2915 4576 3792 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 11054 4604 11060 4616
rect 9263 4576 11060 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 1104 4378 10856 4400
rect 1104 4326 3398 4378
rect 3450 4326 3462 4378
rect 3514 4326 3526 4378
rect 3578 4326 3590 4378
rect 3642 4326 3654 4378
rect 3706 4326 5846 4378
rect 5898 4326 5910 4378
rect 5962 4326 5974 4378
rect 6026 4326 6038 4378
rect 6090 4326 6102 4378
rect 6154 4326 8294 4378
rect 8346 4326 8358 4378
rect 8410 4326 8422 4378
rect 8474 4326 8486 4378
rect 8538 4326 8550 4378
rect 8602 4326 10856 4378
rect 1104 4304 10856 4326
rect 750 3884 756 3936
rect 808 3924 814 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 808 3896 2513 3924
rect 808 3884 814 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 5166 3924 5172 3936
rect 3743 3896 5172 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 6696 3896 7757 3924
rect 6696 3884 6702 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 9033 3927 9091 3933
rect 9033 3924 9045 3927
rect 8168 3896 9045 3924
rect 8168 3884 8174 3896
rect 9033 3893 9045 3896
rect 9079 3893 9091 3927
rect 9033 3887 9091 3893
rect 1104 3834 10856 3856
rect 1104 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 2302 3834
rect 2354 3782 2366 3834
rect 2418 3782 2430 3834
rect 2482 3782 4622 3834
rect 4674 3782 4686 3834
rect 4738 3782 4750 3834
rect 4802 3782 4814 3834
rect 4866 3782 4878 3834
rect 4930 3782 7070 3834
rect 7122 3782 7134 3834
rect 7186 3782 7198 3834
rect 7250 3782 7262 3834
rect 7314 3782 7326 3834
rect 7378 3782 9518 3834
rect 9570 3782 9582 3834
rect 9634 3782 9646 3834
rect 9698 3782 9710 3834
rect 9762 3782 9774 3834
rect 9826 3782 10856 3834
rect 1104 3760 10856 3782
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2556 3488 2697 3516
rect 2556 3476 2562 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9398 3516 9404 3528
rect 9263 3488 9404 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 1104 3290 10856 3312
rect 1104 3238 3398 3290
rect 3450 3238 3462 3290
rect 3514 3238 3526 3290
rect 3578 3238 3590 3290
rect 3642 3238 3654 3290
rect 3706 3238 5846 3290
rect 5898 3238 5910 3290
rect 5962 3238 5974 3290
rect 6026 3238 6038 3290
rect 6090 3238 6102 3290
rect 6154 3238 8294 3290
rect 8346 3238 8358 3290
rect 8410 3238 8422 3290
rect 8474 3238 8486 3290
rect 8538 3238 8550 3290
rect 8602 3238 10856 3290
rect 1104 3216 10856 3238
rect 1104 2746 10856 2768
rect 1104 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 2302 2746
rect 2354 2694 2366 2746
rect 2418 2694 2430 2746
rect 2482 2694 4622 2746
rect 4674 2694 4686 2746
rect 4738 2694 4750 2746
rect 4802 2694 4814 2746
rect 4866 2694 4878 2746
rect 4930 2694 7070 2746
rect 7122 2694 7134 2746
rect 7186 2694 7198 2746
rect 7250 2694 7262 2746
rect 7314 2694 7326 2746
rect 7378 2694 9518 2746
rect 9570 2694 9582 2746
rect 9634 2694 9646 2746
rect 9698 2694 9710 2746
rect 9762 2694 9774 2746
rect 9826 2694 10856 2746
rect 1104 2672 10856 2694
rect 1104 2202 10856 2224
rect 1104 2150 3398 2202
rect 3450 2150 3462 2202
rect 3514 2150 3526 2202
rect 3578 2150 3590 2202
rect 3642 2150 3654 2202
rect 3706 2150 5846 2202
rect 5898 2150 5910 2202
rect 5962 2150 5974 2202
rect 6026 2150 6038 2202
rect 6090 2150 6102 2202
rect 6154 2150 8294 2202
rect 8346 2150 8358 2202
rect 8410 2150 8422 2202
rect 8474 2150 8486 2202
rect 8538 2150 8550 2202
rect 8602 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 2302 11398 2354 11450
rect 2366 11398 2418 11450
rect 2430 11398 2482 11450
rect 4622 11398 4674 11450
rect 4686 11398 4738 11450
rect 4750 11398 4802 11450
rect 4814 11398 4866 11450
rect 4878 11398 4930 11450
rect 7070 11398 7122 11450
rect 7134 11398 7186 11450
rect 7198 11398 7250 11450
rect 7262 11398 7314 11450
rect 7326 11398 7378 11450
rect 9518 11398 9570 11450
rect 9582 11398 9634 11450
rect 9646 11398 9698 11450
rect 9710 11398 9762 11450
rect 9774 11398 9826 11450
rect 3398 10854 3450 10906
rect 3462 10854 3514 10906
rect 3526 10854 3578 10906
rect 3590 10854 3642 10906
rect 3654 10854 3706 10906
rect 5846 10854 5898 10906
rect 5910 10854 5962 10906
rect 5974 10854 6026 10906
rect 6038 10854 6090 10906
rect 6102 10854 6154 10906
rect 8294 10854 8346 10906
rect 8358 10854 8410 10906
rect 8422 10854 8474 10906
rect 8486 10854 8538 10906
rect 8550 10854 8602 10906
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 2302 10310 2354 10362
rect 2366 10310 2418 10362
rect 2430 10310 2482 10362
rect 4622 10310 4674 10362
rect 4686 10310 4738 10362
rect 4750 10310 4802 10362
rect 4814 10310 4866 10362
rect 4878 10310 4930 10362
rect 7070 10310 7122 10362
rect 7134 10310 7186 10362
rect 7198 10310 7250 10362
rect 7262 10310 7314 10362
rect 7326 10310 7378 10362
rect 9518 10310 9570 10362
rect 9582 10310 9634 10362
rect 9646 10310 9698 10362
rect 9710 10310 9762 10362
rect 9774 10310 9826 10362
rect 3398 9766 3450 9818
rect 3462 9766 3514 9818
rect 3526 9766 3578 9818
rect 3590 9766 3642 9818
rect 3654 9766 3706 9818
rect 5846 9766 5898 9818
rect 5910 9766 5962 9818
rect 5974 9766 6026 9818
rect 6038 9766 6090 9818
rect 6102 9766 6154 9818
rect 8294 9766 8346 9818
rect 8358 9766 8410 9818
rect 8422 9766 8474 9818
rect 8486 9766 8538 9818
rect 8550 9766 8602 9818
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 2302 9222 2354 9274
rect 2366 9222 2418 9274
rect 2430 9222 2482 9274
rect 4622 9222 4674 9274
rect 4686 9222 4738 9274
rect 4750 9222 4802 9274
rect 4814 9222 4866 9274
rect 4878 9222 4930 9274
rect 7070 9222 7122 9274
rect 7134 9222 7186 9274
rect 7198 9222 7250 9274
rect 7262 9222 7314 9274
rect 7326 9222 7378 9274
rect 9518 9222 9570 9274
rect 9582 9222 9634 9274
rect 9646 9222 9698 9274
rect 9710 9222 9762 9274
rect 9774 9222 9826 9274
rect 3398 8678 3450 8730
rect 3462 8678 3514 8730
rect 3526 8678 3578 8730
rect 3590 8678 3642 8730
rect 3654 8678 3706 8730
rect 5846 8678 5898 8730
rect 5910 8678 5962 8730
rect 5974 8678 6026 8730
rect 6038 8678 6090 8730
rect 6102 8678 6154 8730
rect 8294 8678 8346 8730
rect 8358 8678 8410 8730
rect 8422 8678 8474 8730
rect 8486 8678 8538 8730
rect 8550 8678 8602 8730
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 2302 8134 2354 8186
rect 2366 8134 2418 8186
rect 2430 8134 2482 8186
rect 4622 8134 4674 8186
rect 4686 8134 4738 8186
rect 4750 8134 4802 8186
rect 4814 8134 4866 8186
rect 4878 8134 4930 8186
rect 7070 8134 7122 8186
rect 7134 8134 7186 8186
rect 7198 8134 7250 8186
rect 7262 8134 7314 8186
rect 7326 8134 7378 8186
rect 9518 8134 9570 8186
rect 9582 8134 9634 8186
rect 9646 8134 9698 8186
rect 9710 8134 9762 8186
rect 9774 8134 9826 8186
rect 3398 7590 3450 7642
rect 3462 7590 3514 7642
rect 3526 7590 3578 7642
rect 3590 7590 3642 7642
rect 3654 7590 3706 7642
rect 5846 7590 5898 7642
rect 5910 7590 5962 7642
rect 5974 7590 6026 7642
rect 6038 7590 6090 7642
rect 6102 7590 6154 7642
rect 8294 7590 8346 7642
rect 8358 7590 8410 7642
rect 8422 7590 8474 7642
rect 8486 7590 8538 7642
rect 8550 7590 8602 7642
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 2302 7046 2354 7098
rect 2366 7046 2418 7098
rect 2430 7046 2482 7098
rect 4622 7046 4674 7098
rect 4686 7046 4738 7098
rect 4750 7046 4802 7098
rect 4814 7046 4866 7098
rect 4878 7046 4930 7098
rect 7070 7046 7122 7098
rect 7134 7046 7186 7098
rect 7198 7046 7250 7098
rect 7262 7046 7314 7098
rect 7326 7046 7378 7098
rect 9518 7046 9570 7098
rect 9582 7046 9634 7098
rect 9646 7046 9698 7098
rect 9710 7046 9762 7098
rect 9774 7046 9826 7098
rect 3398 6502 3450 6554
rect 3462 6502 3514 6554
rect 3526 6502 3578 6554
rect 3590 6502 3642 6554
rect 3654 6502 3706 6554
rect 5846 6502 5898 6554
rect 5910 6502 5962 6554
rect 5974 6502 6026 6554
rect 6038 6502 6090 6554
rect 6102 6502 6154 6554
rect 8294 6502 8346 6554
rect 8358 6502 8410 6554
rect 8422 6502 8474 6554
rect 8486 6502 8538 6554
rect 8550 6502 8602 6554
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 2302 5958 2354 6010
rect 2366 5958 2418 6010
rect 2430 5958 2482 6010
rect 4622 5958 4674 6010
rect 4686 5958 4738 6010
rect 4750 5958 4802 6010
rect 4814 5958 4866 6010
rect 4878 5958 4930 6010
rect 7070 5958 7122 6010
rect 7134 5958 7186 6010
rect 7198 5958 7250 6010
rect 7262 5958 7314 6010
rect 7326 5958 7378 6010
rect 9518 5958 9570 6010
rect 9582 5958 9634 6010
rect 9646 5958 9698 6010
rect 9710 5958 9762 6010
rect 9774 5958 9826 6010
rect 3398 5414 3450 5466
rect 3462 5414 3514 5466
rect 3526 5414 3578 5466
rect 3590 5414 3642 5466
rect 3654 5414 3706 5466
rect 5846 5414 5898 5466
rect 5910 5414 5962 5466
rect 5974 5414 6026 5466
rect 6038 5414 6090 5466
rect 6102 5414 6154 5466
rect 8294 5414 8346 5466
rect 8358 5414 8410 5466
rect 8422 5414 8474 5466
rect 8486 5414 8538 5466
rect 8550 5414 8602 5466
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 2302 4870 2354 4922
rect 2366 4870 2418 4922
rect 2430 4870 2482 4922
rect 4622 4870 4674 4922
rect 4686 4870 4738 4922
rect 4750 4870 4802 4922
rect 4814 4870 4866 4922
rect 4878 4870 4930 4922
rect 7070 4870 7122 4922
rect 7134 4870 7186 4922
rect 7198 4870 7250 4922
rect 7262 4870 7314 4922
rect 7326 4870 7378 4922
rect 9518 4870 9570 4922
rect 9582 4870 9634 4922
rect 9646 4870 9698 4922
rect 9710 4870 9762 4922
rect 9774 4870 9826 4922
rect 3792 4564 3844 4616
rect 11060 4564 11112 4616
rect 3398 4326 3450 4378
rect 3462 4326 3514 4378
rect 3526 4326 3578 4378
rect 3590 4326 3642 4378
rect 3654 4326 3706 4378
rect 5846 4326 5898 4378
rect 5910 4326 5962 4378
rect 5974 4326 6026 4378
rect 6038 4326 6090 4378
rect 6102 4326 6154 4378
rect 8294 4326 8346 4378
rect 8358 4326 8410 4378
rect 8422 4326 8474 4378
rect 8486 4326 8538 4378
rect 8550 4326 8602 4378
rect 756 3884 808 3936
rect 5172 3884 5224 3936
rect 6644 3884 6696 3936
rect 8116 3884 8168 3936
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 2302 3782 2354 3834
rect 2366 3782 2418 3834
rect 2430 3782 2482 3834
rect 4622 3782 4674 3834
rect 4686 3782 4738 3834
rect 4750 3782 4802 3834
rect 4814 3782 4866 3834
rect 4878 3782 4930 3834
rect 7070 3782 7122 3834
rect 7134 3782 7186 3834
rect 7198 3782 7250 3834
rect 7262 3782 7314 3834
rect 7326 3782 7378 3834
rect 9518 3782 9570 3834
rect 9582 3782 9634 3834
rect 9646 3782 9698 3834
rect 9710 3782 9762 3834
rect 9774 3782 9826 3834
rect 2504 3476 2556 3528
rect 9404 3476 9456 3528
rect 3398 3238 3450 3290
rect 3462 3238 3514 3290
rect 3526 3238 3578 3290
rect 3590 3238 3642 3290
rect 3654 3238 3706 3290
rect 5846 3238 5898 3290
rect 5910 3238 5962 3290
rect 5974 3238 6026 3290
rect 6038 3238 6090 3290
rect 6102 3238 6154 3290
rect 8294 3238 8346 3290
rect 8358 3238 8410 3290
rect 8422 3238 8474 3290
rect 8486 3238 8538 3290
rect 8550 3238 8602 3290
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 2302 2694 2354 2746
rect 2366 2694 2418 2746
rect 2430 2694 2482 2746
rect 4622 2694 4674 2746
rect 4686 2694 4738 2746
rect 4750 2694 4802 2746
rect 4814 2694 4866 2746
rect 4878 2694 4930 2746
rect 7070 2694 7122 2746
rect 7134 2694 7186 2746
rect 7198 2694 7250 2746
rect 7262 2694 7314 2746
rect 7326 2694 7378 2746
rect 9518 2694 9570 2746
rect 9582 2694 9634 2746
rect 9646 2694 9698 2746
rect 9710 2694 9762 2746
rect 9774 2694 9826 2746
rect 3398 2150 3450 2202
rect 3462 2150 3514 2202
rect 3526 2150 3578 2202
rect 3590 2150 3642 2202
rect 3654 2150 3706 2202
rect 5846 2150 5898 2202
rect 5910 2150 5962 2202
rect 5974 2150 6026 2202
rect 6038 2150 6090 2202
rect 6102 2150 6154 2202
rect 8294 2150 8346 2202
rect 8358 2150 8410 2202
rect 8422 2150 8474 2202
rect 8486 2150 8538 2202
rect 8550 2150 8602 2202
<< metal2 >>
rect 2174 11452 2482 11461
rect 2174 11450 2180 11452
rect 2236 11450 2260 11452
rect 2316 11450 2340 11452
rect 2396 11450 2420 11452
rect 2476 11450 2482 11452
rect 2236 11398 2238 11450
rect 2418 11398 2420 11450
rect 2174 11396 2180 11398
rect 2236 11396 2260 11398
rect 2316 11396 2340 11398
rect 2396 11396 2420 11398
rect 2476 11396 2482 11398
rect 2174 11387 2482 11396
rect 4622 11452 4930 11461
rect 4622 11450 4628 11452
rect 4684 11450 4708 11452
rect 4764 11450 4788 11452
rect 4844 11450 4868 11452
rect 4924 11450 4930 11452
rect 4684 11398 4686 11450
rect 4866 11398 4868 11450
rect 4622 11396 4628 11398
rect 4684 11396 4708 11398
rect 4764 11396 4788 11398
rect 4844 11396 4868 11398
rect 4924 11396 4930 11398
rect 4622 11387 4930 11396
rect 7070 11452 7378 11461
rect 7070 11450 7076 11452
rect 7132 11450 7156 11452
rect 7212 11450 7236 11452
rect 7292 11450 7316 11452
rect 7372 11450 7378 11452
rect 7132 11398 7134 11450
rect 7314 11398 7316 11450
rect 7070 11396 7076 11398
rect 7132 11396 7156 11398
rect 7212 11396 7236 11398
rect 7292 11396 7316 11398
rect 7372 11396 7378 11398
rect 7070 11387 7378 11396
rect 9518 11452 9826 11461
rect 9518 11450 9524 11452
rect 9580 11450 9604 11452
rect 9660 11450 9684 11452
rect 9740 11450 9764 11452
rect 9820 11450 9826 11452
rect 9580 11398 9582 11450
rect 9762 11398 9764 11450
rect 9518 11396 9524 11398
rect 9580 11396 9604 11398
rect 9660 11396 9684 11398
rect 9740 11396 9764 11398
rect 9820 11396 9826 11398
rect 9518 11387 9826 11396
rect 3398 10908 3706 10917
rect 3398 10906 3404 10908
rect 3460 10906 3484 10908
rect 3540 10906 3564 10908
rect 3620 10906 3644 10908
rect 3700 10906 3706 10908
rect 3460 10854 3462 10906
rect 3642 10854 3644 10906
rect 3398 10852 3404 10854
rect 3460 10852 3484 10854
rect 3540 10852 3564 10854
rect 3620 10852 3644 10854
rect 3700 10852 3706 10854
rect 3398 10843 3706 10852
rect 5846 10908 6154 10917
rect 5846 10906 5852 10908
rect 5908 10906 5932 10908
rect 5988 10906 6012 10908
rect 6068 10906 6092 10908
rect 6148 10906 6154 10908
rect 5908 10854 5910 10906
rect 6090 10854 6092 10906
rect 5846 10852 5852 10854
rect 5908 10852 5932 10854
rect 5988 10852 6012 10854
rect 6068 10852 6092 10854
rect 6148 10852 6154 10854
rect 5846 10843 6154 10852
rect 8294 10908 8602 10917
rect 8294 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8540 10908
rect 8596 10906 8602 10908
rect 8356 10854 8358 10906
rect 8538 10854 8540 10906
rect 8294 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8540 10854
rect 8596 10852 8602 10854
rect 8294 10843 8602 10852
rect 2174 10364 2482 10373
rect 2174 10362 2180 10364
rect 2236 10362 2260 10364
rect 2316 10362 2340 10364
rect 2396 10362 2420 10364
rect 2476 10362 2482 10364
rect 2236 10310 2238 10362
rect 2418 10310 2420 10362
rect 2174 10308 2180 10310
rect 2236 10308 2260 10310
rect 2316 10308 2340 10310
rect 2396 10308 2420 10310
rect 2476 10308 2482 10310
rect 2174 10299 2482 10308
rect 4622 10364 4930 10373
rect 4622 10362 4628 10364
rect 4684 10362 4708 10364
rect 4764 10362 4788 10364
rect 4844 10362 4868 10364
rect 4924 10362 4930 10364
rect 4684 10310 4686 10362
rect 4866 10310 4868 10362
rect 4622 10308 4628 10310
rect 4684 10308 4708 10310
rect 4764 10308 4788 10310
rect 4844 10308 4868 10310
rect 4924 10308 4930 10310
rect 4622 10299 4930 10308
rect 7070 10364 7378 10373
rect 7070 10362 7076 10364
rect 7132 10362 7156 10364
rect 7212 10362 7236 10364
rect 7292 10362 7316 10364
rect 7372 10362 7378 10364
rect 7132 10310 7134 10362
rect 7314 10310 7316 10362
rect 7070 10308 7076 10310
rect 7132 10308 7156 10310
rect 7212 10308 7236 10310
rect 7292 10308 7316 10310
rect 7372 10308 7378 10310
rect 7070 10299 7378 10308
rect 9518 10364 9826 10373
rect 9518 10362 9524 10364
rect 9580 10362 9604 10364
rect 9660 10362 9684 10364
rect 9740 10362 9764 10364
rect 9820 10362 9826 10364
rect 9580 10310 9582 10362
rect 9762 10310 9764 10362
rect 9518 10308 9524 10310
rect 9580 10308 9604 10310
rect 9660 10308 9684 10310
rect 9740 10308 9764 10310
rect 9820 10308 9826 10310
rect 9518 10299 9826 10308
rect 3398 9820 3706 9829
rect 3398 9818 3404 9820
rect 3460 9818 3484 9820
rect 3540 9818 3564 9820
rect 3620 9818 3644 9820
rect 3700 9818 3706 9820
rect 3460 9766 3462 9818
rect 3642 9766 3644 9818
rect 3398 9764 3404 9766
rect 3460 9764 3484 9766
rect 3540 9764 3564 9766
rect 3620 9764 3644 9766
rect 3700 9764 3706 9766
rect 3398 9755 3706 9764
rect 5846 9820 6154 9829
rect 5846 9818 5852 9820
rect 5908 9818 5932 9820
rect 5988 9818 6012 9820
rect 6068 9818 6092 9820
rect 6148 9818 6154 9820
rect 5908 9766 5910 9818
rect 6090 9766 6092 9818
rect 5846 9764 5852 9766
rect 5908 9764 5932 9766
rect 5988 9764 6012 9766
rect 6068 9764 6092 9766
rect 6148 9764 6154 9766
rect 5846 9755 6154 9764
rect 8294 9820 8602 9829
rect 8294 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8540 9820
rect 8596 9818 8602 9820
rect 8356 9766 8358 9818
rect 8538 9766 8540 9818
rect 8294 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8540 9766
rect 8596 9764 8602 9766
rect 8294 9755 8602 9764
rect 2174 9276 2482 9285
rect 2174 9274 2180 9276
rect 2236 9274 2260 9276
rect 2316 9274 2340 9276
rect 2396 9274 2420 9276
rect 2476 9274 2482 9276
rect 2236 9222 2238 9274
rect 2418 9222 2420 9274
rect 2174 9220 2180 9222
rect 2236 9220 2260 9222
rect 2316 9220 2340 9222
rect 2396 9220 2420 9222
rect 2476 9220 2482 9222
rect 2174 9211 2482 9220
rect 4622 9276 4930 9285
rect 4622 9274 4628 9276
rect 4684 9274 4708 9276
rect 4764 9274 4788 9276
rect 4844 9274 4868 9276
rect 4924 9274 4930 9276
rect 4684 9222 4686 9274
rect 4866 9222 4868 9274
rect 4622 9220 4628 9222
rect 4684 9220 4708 9222
rect 4764 9220 4788 9222
rect 4844 9220 4868 9222
rect 4924 9220 4930 9222
rect 4622 9211 4930 9220
rect 7070 9276 7378 9285
rect 7070 9274 7076 9276
rect 7132 9274 7156 9276
rect 7212 9274 7236 9276
rect 7292 9274 7316 9276
rect 7372 9274 7378 9276
rect 7132 9222 7134 9274
rect 7314 9222 7316 9274
rect 7070 9220 7076 9222
rect 7132 9220 7156 9222
rect 7212 9220 7236 9222
rect 7292 9220 7316 9222
rect 7372 9220 7378 9222
rect 7070 9211 7378 9220
rect 9518 9276 9826 9285
rect 9518 9274 9524 9276
rect 9580 9274 9604 9276
rect 9660 9274 9684 9276
rect 9740 9274 9764 9276
rect 9820 9274 9826 9276
rect 9580 9222 9582 9274
rect 9762 9222 9764 9274
rect 9518 9220 9524 9222
rect 9580 9220 9604 9222
rect 9660 9220 9684 9222
rect 9740 9220 9764 9222
rect 9820 9220 9826 9222
rect 9518 9211 9826 9220
rect 3398 8732 3706 8741
rect 3398 8730 3404 8732
rect 3460 8730 3484 8732
rect 3540 8730 3564 8732
rect 3620 8730 3644 8732
rect 3700 8730 3706 8732
rect 3460 8678 3462 8730
rect 3642 8678 3644 8730
rect 3398 8676 3404 8678
rect 3460 8676 3484 8678
rect 3540 8676 3564 8678
rect 3620 8676 3644 8678
rect 3700 8676 3706 8678
rect 3398 8667 3706 8676
rect 5846 8732 6154 8741
rect 5846 8730 5852 8732
rect 5908 8730 5932 8732
rect 5988 8730 6012 8732
rect 6068 8730 6092 8732
rect 6148 8730 6154 8732
rect 5908 8678 5910 8730
rect 6090 8678 6092 8730
rect 5846 8676 5852 8678
rect 5908 8676 5932 8678
rect 5988 8676 6012 8678
rect 6068 8676 6092 8678
rect 6148 8676 6154 8678
rect 5846 8667 6154 8676
rect 8294 8732 8602 8741
rect 8294 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8540 8732
rect 8596 8730 8602 8732
rect 8356 8678 8358 8730
rect 8538 8678 8540 8730
rect 8294 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8540 8678
rect 8596 8676 8602 8678
rect 8294 8667 8602 8676
rect 2174 8188 2482 8197
rect 2174 8186 2180 8188
rect 2236 8186 2260 8188
rect 2316 8186 2340 8188
rect 2396 8186 2420 8188
rect 2476 8186 2482 8188
rect 2236 8134 2238 8186
rect 2418 8134 2420 8186
rect 2174 8132 2180 8134
rect 2236 8132 2260 8134
rect 2316 8132 2340 8134
rect 2396 8132 2420 8134
rect 2476 8132 2482 8134
rect 2174 8123 2482 8132
rect 4622 8188 4930 8197
rect 4622 8186 4628 8188
rect 4684 8186 4708 8188
rect 4764 8186 4788 8188
rect 4844 8186 4868 8188
rect 4924 8186 4930 8188
rect 4684 8134 4686 8186
rect 4866 8134 4868 8186
rect 4622 8132 4628 8134
rect 4684 8132 4708 8134
rect 4764 8132 4788 8134
rect 4844 8132 4868 8134
rect 4924 8132 4930 8134
rect 4622 8123 4930 8132
rect 7070 8188 7378 8197
rect 7070 8186 7076 8188
rect 7132 8186 7156 8188
rect 7212 8186 7236 8188
rect 7292 8186 7316 8188
rect 7372 8186 7378 8188
rect 7132 8134 7134 8186
rect 7314 8134 7316 8186
rect 7070 8132 7076 8134
rect 7132 8132 7156 8134
rect 7212 8132 7236 8134
rect 7292 8132 7316 8134
rect 7372 8132 7378 8134
rect 7070 8123 7378 8132
rect 9518 8188 9826 8197
rect 9518 8186 9524 8188
rect 9580 8186 9604 8188
rect 9660 8186 9684 8188
rect 9740 8186 9764 8188
rect 9820 8186 9826 8188
rect 9580 8134 9582 8186
rect 9762 8134 9764 8186
rect 9518 8132 9524 8134
rect 9580 8132 9604 8134
rect 9660 8132 9684 8134
rect 9740 8132 9764 8134
rect 9820 8132 9826 8134
rect 9518 8123 9826 8132
rect 3398 7644 3706 7653
rect 3398 7642 3404 7644
rect 3460 7642 3484 7644
rect 3540 7642 3564 7644
rect 3620 7642 3644 7644
rect 3700 7642 3706 7644
rect 3460 7590 3462 7642
rect 3642 7590 3644 7642
rect 3398 7588 3404 7590
rect 3460 7588 3484 7590
rect 3540 7588 3564 7590
rect 3620 7588 3644 7590
rect 3700 7588 3706 7590
rect 3398 7579 3706 7588
rect 5846 7644 6154 7653
rect 5846 7642 5852 7644
rect 5908 7642 5932 7644
rect 5988 7642 6012 7644
rect 6068 7642 6092 7644
rect 6148 7642 6154 7644
rect 5908 7590 5910 7642
rect 6090 7590 6092 7642
rect 5846 7588 5852 7590
rect 5908 7588 5932 7590
rect 5988 7588 6012 7590
rect 6068 7588 6092 7590
rect 6148 7588 6154 7590
rect 5846 7579 6154 7588
rect 8294 7644 8602 7653
rect 8294 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8540 7644
rect 8596 7642 8602 7644
rect 8356 7590 8358 7642
rect 8538 7590 8540 7642
rect 8294 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8540 7590
rect 8596 7588 8602 7590
rect 8294 7579 8602 7588
rect 2174 7100 2482 7109
rect 2174 7098 2180 7100
rect 2236 7098 2260 7100
rect 2316 7098 2340 7100
rect 2396 7098 2420 7100
rect 2476 7098 2482 7100
rect 2236 7046 2238 7098
rect 2418 7046 2420 7098
rect 2174 7044 2180 7046
rect 2236 7044 2260 7046
rect 2316 7044 2340 7046
rect 2396 7044 2420 7046
rect 2476 7044 2482 7046
rect 2174 7035 2482 7044
rect 4622 7100 4930 7109
rect 4622 7098 4628 7100
rect 4684 7098 4708 7100
rect 4764 7098 4788 7100
rect 4844 7098 4868 7100
rect 4924 7098 4930 7100
rect 4684 7046 4686 7098
rect 4866 7046 4868 7098
rect 4622 7044 4628 7046
rect 4684 7044 4708 7046
rect 4764 7044 4788 7046
rect 4844 7044 4868 7046
rect 4924 7044 4930 7046
rect 4622 7035 4930 7044
rect 7070 7100 7378 7109
rect 7070 7098 7076 7100
rect 7132 7098 7156 7100
rect 7212 7098 7236 7100
rect 7292 7098 7316 7100
rect 7372 7098 7378 7100
rect 7132 7046 7134 7098
rect 7314 7046 7316 7098
rect 7070 7044 7076 7046
rect 7132 7044 7156 7046
rect 7212 7044 7236 7046
rect 7292 7044 7316 7046
rect 7372 7044 7378 7046
rect 7070 7035 7378 7044
rect 9518 7100 9826 7109
rect 9518 7098 9524 7100
rect 9580 7098 9604 7100
rect 9660 7098 9684 7100
rect 9740 7098 9764 7100
rect 9820 7098 9826 7100
rect 9580 7046 9582 7098
rect 9762 7046 9764 7098
rect 9518 7044 9524 7046
rect 9580 7044 9604 7046
rect 9660 7044 9684 7046
rect 9740 7044 9764 7046
rect 9820 7044 9826 7046
rect 9518 7035 9826 7044
rect 3398 6556 3706 6565
rect 3398 6554 3404 6556
rect 3460 6554 3484 6556
rect 3540 6554 3564 6556
rect 3620 6554 3644 6556
rect 3700 6554 3706 6556
rect 3460 6502 3462 6554
rect 3642 6502 3644 6554
rect 3398 6500 3404 6502
rect 3460 6500 3484 6502
rect 3540 6500 3564 6502
rect 3620 6500 3644 6502
rect 3700 6500 3706 6502
rect 3398 6491 3706 6500
rect 5846 6556 6154 6565
rect 5846 6554 5852 6556
rect 5908 6554 5932 6556
rect 5988 6554 6012 6556
rect 6068 6554 6092 6556
rect 6148 6554 6154 6556
rect 5908 6502 5910 6554
rect 6090 6502 6092 6554
rect 5846 6500 5852 6502
rect 5908 6500 5932 6502
rect 5988 6500 6012 6502
rect 6068 6500 6092 6502
rect 6148 6500 6154 6502
rect 5846 6491 6154 6500
rect 8294 6556 8602 6565
rect 8294 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8540 6556
rect 8596 6554 8602 6556
rect 8356 6502 8358 6554
rect 8538 6502 8540 6554
rect 8294 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8540 6502
rect 8596 6500 8602 6502
rect 8294 6491 8602 6500
rect 2174 6012 2482 6021
rect 2174 6010 2180 6012
rect 2236 6010 2260 6012
rect 2316 6010 2340 6012
rect 2396 6010 2420 6012
rect 2476 6010 2482 6012
rect 2236 5958 2238 6010
rect 2418 5958 2420 6010
rect 2174 5956 2180 5958
rect 2236 5956 2260 5958
rect 2316 5956 2340 5958
rect 2396 5956 2420 5958
rect 2476 5956 2482 5958
rect 2174 5947 2482 5956
rect 4622 6012 4930 6021
rect 4622 6010 4628 6012
rect 4684 6010 4708 6012
rect 4764 6010 4788 6012
rect 4844 6010 4868 6012
rect 4924 6010 4930 6012
rect 4684 5958 4686 6010
rect 4866 5958 4868 6010
rect 4622 5956 4628 5958
rect 4684 5956 4708 5958
rect 4764 5956 4788 5958
rect 4844 5956 4868 5958
rect 4924 5956 4930 5958
rect 4622 5947 4930 5956
rect 7070 6012 7378 6021
rect 7070 6010 7076 6012
rect 7132 6010 7156 6012
rect 7212 6010 7236 6012
rect 7292 6010 7316 6012
rect 7372 6010 7378 6012
rect 7132 5958 7134 6010
rect 7314 5958 7316 6010
rect 7070 5956 7076 5958
rect 7132 5956 7156 5958
rect 7212 5956 7236 5958
rect 7292 5956 7316 5958
rect 7372 5956 7378 5958
rect 7070 5947 7378 5956
rect 9518 6012 9826 6021
rect 9518 6010 9524 6012
rect 9580 6010 9604 6012
rect 9660 6010 9684 6012
rect 9740 6010 9764 6012
rect 9820 6010 9826 6012
rect 9580 5958 9582 6010
rect 9762 5958 9764 6010
rect 9518 5956 9524 5958
rect 9580 5956 9604 5958
rect 9660 5956 9684 5958
rect 9740 5956 9764 5958
rect 9820 5956 9826 5958
rect 9518 5947 9826 5956
rect 3398 5468 3706 5477
rect 3398 5466 3404 5468
rect 3460 5466 3484 5468
rect 3540 5466 3564 5468
rect 3620 5466 3644 5468
rect 3700 5466 3706 5468
rect 3460 5414 3462 5466
rect 3642 5414 3644 5466
rect 3398 5412 3404 5414
rect 3460 5412 3484 5414
rect 3540 5412 3564 5414
rect 3620 5412 3644 5414
rect 3700 5412 3706 5414
rect 3398 5403 3706 5412
rect 5846 5468 6154 5477
rect 5846 5466 5852 5468
rect 5908 5466 5932 5468
rect 5988 5466 6012 5468
rect 6068 5466 6092 5468
rect 6148 5466 6154 5468
rect 5908 5414 5910 5466
rect 6090 5414 6092 5466
rect 5846 5412 5852 5414
rect 5908 5412 5932 5414
rect 5988 5412 6012 5414
rect 6068 5412 6092 5414
rect 6148 5412 6154 5414
rect 5846 5403 6154 5412
rect 8294 5468 8602 5477
rect 8294 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8540 5468
rect 8596 5466 8602 5468
rect 8356 5414 8358 5466
rect 8538 5414 8540 5466
rect 8294 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8540 5414
rect 8596 5412 8602 5414
rect 8294 5403 8602 5412
rect 2174 4924 2482 4933
rect 2174 4922 2180 4924
rect 2236 4922 2260 4924
rect 2316 4922 2340 4924
rect 2396 4922 2420 4924
rect 2476 4922 2482 4924
rect 2236 4870 2238 4922
rect 2418 4870 2420 4922
rect 2174 4868 2180 4870
rect 2236 4868 2260 4870
rect 2316 4868 2340 4870
rect 2396 4868 2420 4870
rect 2476 4868 2482 4870
rect 2174 4859 2482 4868
rect 4622 4924 4930 4933
rect 4622 4922 4628 4924
rect 4684 4922 4708 4924
rect 4764 4922 4788 4924
rect 4844 4922 4868 4924
rect 4924 4922 4930 4924
rect 4684 4870 4686 4922
rect 4866 4870 4868 4922
rect 4622 4868 4628 4870
rect 4684 4868 4708 4870
rect 4764 4868 4788 4870
rect 4844 4868 4868 4870
rect 4924 4868 4930 4870
rect 4622 4859 4930 4868
rect 7070 4924 7378 4933
rect 7070 4922 7076 4924
rect 7132 4922 7156 4924
rect 7212 4922 7236 4924
rect 7292 4922 7316 4924
rect 7372 4922 7378 4924
rect 7132 4870 7134 4922
rect 7314 4870 7316 4922
rect 7070 4868 7076 4870
rect 7132 4868 7156 4870
rect 7212 4868 7236 4870
rect 7292 4868 7316 4870
rect 7372 4868 7378 4870
rect 7070 4859 7378 4868
rect 9518 4924 9826 4933
rect 9518 4922 9524 4924
rect 9580 4922 9604 4924
rect 9660 4922 9684 4924
rect 9740 4922 9764 4924
rect 9820 4922 9826 4924
rect 9580 4870 9582 4922
rect 9762 4870 9764 4922
rect 9518 4868 9524 4870
rect 9580 4868 9604 4870
rect 9660 4868 9684 4870
rect 9740 4868 9764 4870
rect 9820 4868 9826 4870
rect 9518 4859 9826 4868
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 3398 4380 3706 4389
rect 3398 4378 3404 4380
rect 3460 4378 3484 4380
rect 3540 4378 3564 4380
rect 3620 4378 3644 4380
rect 3700 4378 3706 4380
rect 3460 4326 3462 4378
rect 3642 4326 3644 4378
rect 3398 4324 3404 4326
rect 3460 4324 3484 4326
rect 3540 4324 3564 4326
rect 3620 4324 3644 4326
rect 3700 4324 3706 4326
rect 3398 4315 3706 4324
rect 756 3936 808 3942
rect 756 3878 808 3884
rect 768 800 796 3878
rect 2174 3836 2482 3845
rect 2174 3834 2180 3836
rect 2236 3834 2260 3836
rect 2316 3834 2340 3836
rect 2396 3834 2420 3836
rect 2476 3834 2482 3836
rect 2236 3782 2238 3834
rect 2418 3782 2420 3834
rect 2174 3780 2180 3782
rect 2236 3780 2260 3782
rect 2316 3780 2340 3782
rect 2396 3780 2420 3782
rect 2476 3780 2482 3782
rect 2174 3771 2482 3780
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2174 2748 2482 2757
rect 2174 2746 2180 2748
rect 2236 2746 2260 2748
rect 2316 2746 2340 2748
rect 2396 2746 2420 2748
rect 2476 2746 2482 2748
rect 2236 2694 2238 2746
rect 2418 2694 2420 2746
rect 2174 2692 2180 2694
rect 2236 2692 2260 2694
rect 2316 2692 2340 2694
rect 2396 2692 2420 2694
rect 2476 2692 2482 2694
rect 2174 2683 2482 2692
rect 2240 870 2360 898
rect 2240 800 2268 870
rect 754 0 810 800
rect 2226 0 2282 800
rect 2332 762 2360 870
rect 2516 762 2544 3470
rect 3398 3292 3706 3301
rect 3398 3290 3404 3292
rect 3460 3290 3484 3292
rect 3540 3290 3564 3292
rect 3620 3290 3644 3292
rect 3700 3290 3706 3292
rect 3460 3238 3462 3290
rect 3642 3238 3644 3290
rect 3398 3236 3404 3238
rect 3460 3236 3484 3238
rect 3540 3236 3564 3238
rect 3620 3236 3644 3238
rect 3700 3236 3706 3238
rect 3398 3227 3706 3236
rect 3398 2204 3706 2213
rect 3398 2202 3404 2204
rect 3460 2202 3484 2204
rect 3540 2202 3564 2204
rect 3620 2202 3644 2204
rect 3700 2202 3706 2204
rect 3460 2150 3462 2202
rect 3642 2150 3644 2202
rect 3398 2148 3404 2150
rect 3460 2148 3484 2150
rect 3540 2148 3564 2150
rect 3620 2148 3644 2150
rect 3700 2148 3706 2150
rect 3398 2139 3706 2148
rect 3804 1986 3832 4558
rect 5846 4380 6154 4389
rect 5846 4378 5852 4380
rect 5908 4378 5932 4380
rect 5988 4378 6012 4380
rect 6068 4378 6092 4380
rect 6148 4378 6154 4380
rect 5908 4326 5910 4378
rect 6090 4326 6092 4378
rect 5846 4324 5852 4326
rect 5908 4324 5932 4326
rect 5988 4324 6012 4326
rect 6068 4324 6092 4326
rect 6148 4324 6154 4326
rect 5846 4315 6154 4324
rect 8294 4380 8602 4389
rect 8294 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8540 4380
rect 8596 4378 8602 4380
rect 8356 4326 8358 4378
rect 8538 4326 8540 4378
rect 8294 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8540 4326
rect 8596 4324 8602 4326
rect 8294 4315 8602 4324
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 4622 3836 4930 3845
rect 4622 3834 4628 3836
rect 4684 3834 4708 3836
rect 4764 3834 4788 3836
rect 4844 3834 4868 3836
rect 4924 3834 4930 3836
rect 4684 3782 4686 3834
rect 4866 3782 4868 3834
rect 4622 3780 4628 3782
rect 4684 3780 4708 3782
rect 4764 3780 4788 3782
rect 4844 3780 4868 3782
rect 4924 3780 4930 3782
rect 4622 3771 4930 3780
rect 4622 2748 4930 2757
rect 4622 2746 4628 2748
rect 4684 2746 4708 2748
rect 4764 2746 4788 2748
rect 4844 2746 4868 2748
rect 4924 2746 4930 2748
rect 4684 2694 4686 2746
rect 4866 2694 4868 2746
rect 4622 2692 4628 2694
rect 4684 2692 4708 2694
rect 4764 2692 4788 2694
rect 4844 2692 4868 2694
rect 4924 2692 4930 2694
rect 4622 2683 4930 2692
rect 3712 1958 3832 1986
rect 3712 800 3740 1958
rect 5184 800 5212 3878
rect 5846 3292 6154 3301
rect 5846 3290 5852 3292
rect 5908 3290 5932 3292
rect 5988 3290 6012 3292
rect 6068 3290 6092 3292
rect 6148 3290 6154 3292
rect 5908 3238 5910 3290
rect 6090 3238 6092 3290
rect 5846 3236 5852 3238
rect 5908 3236 5932 3238
rect 5988 3236 6012 3238
rect 6068 3236 6092 3238
rect 6148 3236 6154 3238
rect 5846 3227 6154 3236
rect 5846 2204 6154 2213
rect 5846 2202 5852 2204
rect 5908 2202 5932 2204
rect 5988 2202 6012 2204
rect 6068 2202 6092 2204
rect 6148 2202 6154 2204
rect 5908 2150 5910 2202
rect 6090 2150 6092 2202
rect 5846 2148 5852 2150
rect 5908 2148 5932 2150
rect 5988 2148 6012 2150
rect 6068 2148 6092 2150
rect 6148 2148 6154 2150
rect 5846 2139 6154 2148
rect 6656 800 6684 3878
rect 7070 3836 7378 3845
rect 7070 3834 7076 3836
rect 7132 3834 7156 3836
rect 7212 3834 7236 3836
rect 7292 3834 7316 3836
rect 7372 3834 7378 3836
rect 7132 3782 7134 3834
rect 7314 3782 7316 3834
rect 7070 3780 7076 3782
rect 7132 3780 7156 3782
rect 7212 3780 7236 3782
rect 7292 3780 7316 3782
rect 7372 3780 7378 3782
rect 7070 3771 7378 3780
rect 7070 2748 7378 2757
rect 7070 2746 7076 2748
rect 7132 2746 7156 2748
rect 7212 2746 7236 2748
rect 7292 2746 7316 2748
rect 7372 2746 7378 2748
rect 7132 2694 7134 2746
rect 7314 2694 7316 2746
rect 7070 2692 7076 2694
rect 7132 2692 7156 2694
rect 7212 2692 7236 2694
rect 7292 2692 7316 2694
rect 7372 2692 7378 2694
rect 7070 2683 7378 2692
rect 8128 800 8156 3878
rect 9518 3836 9826 3845
rect 9518 3834 9524 3836
rect 9580 3834 9604 3836
rect 9660 3834 9684 3836
rect 9740 3834 9764 3836
rect 9820 3834 9826 3836
rect 9580 3782 9582 3834
rect 9762 3782 9764 3834
rect 9518 3780 9524 3782
rect 9580 3780 9604 3782
rect 9660 3780 9684 3782
rect 9740 3780 9764 3782
rect 9820 3780 9826 3782
rect 9518 3771 9826 3780
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8294 3292 8602 3301
rect 8294 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8540 3292
rect 8596 3290 8602 3292
rect 8356 3238 8358 3290
rect 8538 3238 8540 3290
rect 8294 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8540 3238
rect 8596 3236 8602 3238
rect 8294 3227 8602 3236
rect 8294 2204 8602 2213
rect 8294 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8540 2204
rect 8596 2202 8602 2204
rect 8356 2150 8358 2202
rect 8538 2150 8540 2202
rect 8294 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8540 2150
rect 8596 2148 8602 2150
rect 8294 2139 8602 2148
rect 9416 1850 9444 3470
rect 9518 2748 9826 2757
rect 9518 2746 9524 2748
rect 9580 2746 9604 2748
rect 9660 2746 9684 2748
rect 9740 2746 9764 2748
rect 9820 2746 9826 2748
rect 9580 2694 9582 2746
rect 9762 2694 9764 2746
rect 9518 2692 9524 2694
rect 9580 2692 9604 2694
rect 9660 2692 9684 2694
rect 9740 2692 9764 2694
rect 9820 2692 9826 2694
rect 9518 2683 9826 2692
rect 9416 1822 9628 1850
rect 9600 800 9628 1822
rect 11072 800 11100 4558
rect 2332 734 2544 762
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9586 0 9642 800
rect 11058 0 11114 800
<< via2 >>
rect 2180 11450 2236 11452
rect 2260 11450 2316 11452
rect 2340 11450 2396 11452
rect 2420 11450 2476 11452
rect 2180 11398 2226 11450
rect 2226 11398 2236 11450
rect 2260 11398 2290 11450
rect 2290 11398 2302 11450
rect 2302 11398 2316 11450
rect 2340 11398 2354 11450
rect 2354 11398 2366 11450
rect 2366 11398 2396 11450
rect 2420 11398 2430 11450
rect 2430 11398 2476 11450
rect 2180 11396 2236 11398
rect 2260 11396 2316 11398
rect 2340 11396 2396 11398
rect 2420 11396 2476 11398
rect 4628 11450 4684 11452
rect 4708 11450 4764 11452
rect 4788 11450 4844 11452
rect 4868 11450 4924 11452
rect 4628 11398 4674 11450
rect 4674 11398 4684 11450
rect 4708 11398 4738 11450
rect 4738 11398 4750 11450
rect 4750 11398 4764 11450
rect 4788 11398 4802 11450
rect 4802 11398 4814 11450
rect 4814 11398 4844 11450
rect 4868 11398 4878 11450
rect 4878 11398 4924 11450
rect 4628 11396 4684 11398
rect 4708 11396 4764 11398
rect 4788 11396 4844 11398
rect 4868 11396 4924 11398
rect 7076 11450 7132 11452
rect 7156 11450 7212 11452
rect 7236 11450 7292 11452
rect 7316 11450 7372 11452
rect 7076 11398 7122 11450
rect 7122 11398 7132 11450
rect 7156 11398 7186 11450
rect 7186 11398 7198 11450
rect 7198 11398 7212 11450
rect 7236 11398 7250 11450
rect 7250 11398 7262 11450
rect 7262 11398 7292 11450
rect 7316 11398 7326 11450
rect 7326 11398 7372 11450
rect 7076 11396 7132 11398
rect 7156 11396 7212 11398
rect 7236 11396 7292 11398
rect 7316 11396 7372 11398
rect 9524 11450 9580 11452
rect 9604 11450 9660 11452
rect 9684 11450 9740 11452
rect 9764 11450 9820 11452
rect 9524 11398 9570 11450
rect 9570 11398 9580 11450
rect 9604 11398 9634 11450
rect 9634 11398 9646 11450
rect 9646 11398 9660 11450
rect 9684 11398 9698 11450
rect 9698 11398 9710 11450
rect 9710 11398 9740 11450
rect 9764 11398 9774 11450
rect 9774 11398 9820 11450
rect 9524 11396 9580 11398
rect 9604 11396 9660 11398
rect 9684 11396 9740 11398
rect 9764 11396 9820 11398
rect 3404 10906 3460 10908
rect 3484 10906 3540 10908
rect 3564 10906 3620 10908
rect 3644 10906 3700 10908
rect 3404 10854 3450 10906
rect 3450 10854 3460 10906
rect 3484 10854 3514 10906
rect 3514 10854 3526 10906
rect 3526 10854 3540 10906
rect 3564 10854 3578 10906
rect 3578 10854 3590 10906
rect 3590 10854 3620 10906
rect 3644 10854 3654 10906
rect 3654 10854 3700 10906
rect 3404 10852 3460 10854
rect 3484 10852 3540 10854
rect 3564 10852 3620 10854
rect 3644 10852 3700 10854
rect 5852 10906 5908 10908
rect 5932 10906 5988 10908
rect 6012 10906 6068 10908
rect 6092 10906 6148 10908
rect 5852 10854 5898 10906
rect 5898 10854 5908 10906
rect 5932 10854 5962 10906
rect 5962 10854 5974 10906
rect 5974 10854 5988 10906
rect 6012 10854 6026 10906
rect 6026 10854 6038 10906
rect 6038 10854 6068 10906
rect 6092 10854 6102 10906
rect 6102 10854 6148 10906
rect 5852 10852 5908 10854
rect 5932 10852 5988 10854
rect 6012 10852 6068 10854
rect 6092 10852 6148 10854
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8540 10906 8596 10908
rect 8300 10854 8346 10906
rect 8346 10854 8356 10906
rect 8380 10854 8410 10906
rect 8410 10854 8422 10906
rect 8422 10854 8436 10906
rect 8460 10854 8474 10906
rect 8474 10854 8486 10906
rect 8486 10854 8516 10906
rect 8540 10854 8550 10906
rect 8550 10854 8596 10906
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8540 10852 8596 10854
rect 2180 10362 2236 10364
rect 2260 10362 2316 10364
rect 2340 10362 2396 10364
rect 2420 10362 2476 10364
rect 2180 10310 2226 10362
rect 2226 10310 2236 10362
rect 2260 10310 2290 10362
rect 2290 10310 2302 10362
rect 2302 10310 2316 10362
rect 2340 10310 2354 10362
rect 2354 10310 2366 10362
rect 2366 10310 2396 10362
rect 2420 10310 2430 10362
rect 2430 10310 2476 10362
rect 2180 10308 2236 10310
rect 2260 10308 2316 10310
rect 2340 10308 2396 10310
rect 2420 10308 2476 10310
rect 4628 10362 4684 10364
rect 4708 10362 4764 10364
rect 4788 10362 4844 10364
rect 4868 10362 4924 10364
rect 4628 10310 4674 10362
rect 4674 10310 4684 10362
rect 4708 10310 4738 10362
rect 4738 10310 4750 10362
rect 4750 10310 4764 10362
rect 4788 10310 4802 10362
rect 4802 10310 4814 10362
rect 4814 10310 4844 10362
rect 4868 10310 4878 10362
rect 4878 10310 4924 10362
rect 4628 10308 4684 10310
rect 4708 10308 4764 10310
rect 4788 10308 4844 10310
rect 4868 10308 4924 10310
rect 7076 10362 7132 10364
rect 7156 10362 7212 10364
rect 7236 10362 7292 10364
rect 7316 10362 7372 10364
rect 7076 10310 7122 10362
rect 7122 10310 7132 10362
rect 7156 10310 7186 10362
rect 7186 10310 7198 10362
rect 7198 10310 7212 10362
rect 7236 10310 7250 10362
rect 7250 10310 7262 10362
rect 7262 10310 7292 10362
rect 7316 10310 7326 10362
rect 7326 10310 7372 10362
rect 7076 10308 7132 10310
rect 7156 10308 7212 10310
rect 7236 10308 7292 10310
rect 7316 10308 7372 10310
rect 9524 10362 9580 10364
rect 9604 10362 9660 10364
rect 9684 10362 9740 10364
rect 9764 10362 9820 10364
rect 9524 10310 9570 10362
rect 9570 10310 9580 10362
rect 9604 10310 9634 10362
rect 9634 10310 9646 10362
rect 9646 10310 9660 10362
rect 9684 10310 9698 10362
rect 9698 10310 9710 10362
rect 9710 10310 9740 10362
rect 9764 10310 9774 10362
rect 9774 10310 9820 10362
rect 9524 10308 9580 10310
rect 9604 10308 9660 10310
rect 9684 10308 9740 10310
rect 9764 10308 9820 10310
rect 3404 9818 3460 9820
rect 3484 9818 3540 9820
rect 3564 9818 3620 9820
rect 3644 9818 3700 9820
rect 3404 9766 3450 9818
rect 3450 9766 3460 9818
rect 3484 9766 3514 9818
rect 3514 9766 3526 9818
rect 3526 9766 3540 9818
rect 3564 9766 3578 9818
rect 3578 9766 3590 9818
rect 3590 9766 3620 9818
rect 3644 9766 3654 9818
rect 3654 9766 3700 9818
rect 3404 9764 3460 9766
rect 3484 9764 3540 9766
rect 3564 9764 3620 9766
rect 3644 9764 3700 9766
rect 5852 9818 5908 9820
rect 5932 9818 5988 9820
rect 6012 9818 6068 9820
rect 6092 9818 6148 9820
rect 5852 9766 5898 9818
rect 5898 9766 5908 9818
rect 5932 9766 5962 9818
rect 5962 9766 5974 9818
rect 5974 9766 5988 9818
rect 6012 9766 6026 9818
rect 6026 9766 6038 9818
rect 6038 9766 6068 9818
rect 6092 9766 6102 9818
rect 6102 9766 6148 9818
rect 5852 9764 5908 9766
rect 5932 9764 5988 9766
rect 6012 9764 6068 9766
rect 6092 9764 6148 9766
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8540 9818 8596 9820
rect 8300 9766 8346 9818
rect 8346 9766 8356 9818
rect 8380 9766 8410 9818
rect 8410 9766 8422 9818
rect 8422 9766 8436 9818
rect 8460 9766 8474 9818
rect 8474 9766 8486 9818
rect 8486 9766 8516 9818
rect 8540 9766 8550 9818
rect 8550 9766 8596 9818
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8540 9764 8596 9766
rect 2180 9274 2236 9276
rect 2260 9274 2316 9276
rect 2340 9274 2396 9276
rect 2420 9274 2476 9276
rect 2180 9222 2226 9274
rect 2226 9222 2236 9274
rect 2260 9222 2290 9274
rect 2290 9222 2302 9274
rect 2302 9222 2316 9274
rect 2340 9222 2354 9274
rect 2354 9222 2366 9274
rect 2366 9222 2396 9274
rect 2420 9222 2430 9274
rect 2430 9222 2476 9274
rect 2180 9220 2236 9222
rect 2260 9220 2316 9222
rect 2340 9220 2396 9222
rect 2420 9220 2476 9222
rect 4628 9274 4684 9276
rect 4708 9274 4764 9276
rect 4788 9274 4844 9276
rect 4868 9274 4924 9276
rect 4628 9222 4674 9274
rect 4674 9222 4684 9274
rect 4708 9222 4738 9274
rect 4738 9222 4750 9274
rect 4750 9222 4764 9274
rect 4788 9222 4802 9274
rect 4802 9222 4814 9274
rect 4814 9222 4844 9274
rect 4868 9222 4878 9274
rect 4878 9222 4924 9274
rect 4628 9220 4684 9222
rect 4708 9220 4764 9222
rect 4788 9220 4844 9222
rect 4868 9220 4924 9222
rect 7076 9274 7132 9276
rect 7156 9274 7212 9276
rect 7236 9274 7292 9276
rect 7316 9274 7372 9276
rect 7076 9222 7122 9274
rect 7122 9222 7132 9274
rect 7156 9222 7186 9274
rect 7186 9222 7198 9274
rect 7198 9222 7212 9274
rect 7236 9222 7250 9274
rect 7250 9222 7262 9274
rect 7262 9222 7292 9274
rect 7316 9222 7326 9274
rect 7326 9222 7372 9274
rect 7076 9220 7132 9222
rect 7156 9220 7212 9222
rect 7236 9220 7292 9222
rect 7316 9220 7372 9222
rect 9524 9274 9580 9276
rect 9604 9274 9660 9276
rect 9684 9274 9740 9276
rect 9764 9274 9820 9276
rect 9524 9222 9570 9274
rect 9570 9222 9580 9274
rect 9604 9222 9634 9274
rect 9634 9222 9646 9274
rect 9646 9222 9660 9274
rect 9684 9222 9698 9274
rect 9698 9222 9710 9274
rect 9710 9222 9740 9274
rect 9764 9222 9774 9274
rect 9774 9222 9820 9274
rect 9524 9220 9580 9222
rect 9604 9220 9660 9222
rect 9684 9220 9740 9222
rect 9764 9220 9820 9222
rect 3404 8730 3460 8732
rect 3484 8730 3540 8732
rect 3564 8730 3620 8732
rect 3644 8730 3700 8732
rect 3404 8678 3450 8730
rect 3450 8678 3460 8730
rect 3484 8678 3514 8730
rect 3514 8678 3526 8730
rect 3526 8678 3540 8730
rect 3564 8678 3578 8730
rect 3578 8678 3590 8730
rect 3590 8678 3620 8730
rect 3644 8678 3654 8730
rect 3654 8678 3700 8730
rect 3404 8676 3460 8678
rect 3484 8676 3540 8678
rect 3564 8676 3620 8678
rect 3644 8676 3700 8678
rect 5852 8730 5908 8732
rect 5932 8730 5988 8732
rect 6012 8730 6068 8732
rect 6092 8730 6148 8732
rect 5852 8678 5898 8730
rect 5898 8678 5908 8730
rect 5932 8678 5962 8730
rect 5962 8678 5974 8730
rect 5974 8678 5988 8730
rect 6012 8678 6026 8730
rect 6026 8678 6038 8730
rect 6038 8678 6068 8730
rect 6092 8678 6102 8730
rect 6102 8678 6148 8730
rect 5852 8676 5908 8678
rect 5932 8676 5988 8678
rect 6012 8676 6068 8678
rect 6092 8676 6148 8678
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8540 8730 8596 8732
rect 8300 8678 8346 8730
rect 8346 8678 8356 8730
rect 8380 8678 8410 8730
rect 8410 8678 8422 8730
rect 8422 8678 8436 8730
rect 8460 8678 8474 8730
rect 8474 8678 8486 8730
rect 8486 8678 8516 8730
rect 8540 8678 8550 8730
rect 8550 8678 8596 8730
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8540 8676 8596 8678
rect 2180 8186 2236 8188
rect 2260 8186 2316 8188
rect 2340 8186 2396 8188
rect 2420 8186 2476 8188
rect 2180 8134 2226 8186
rect 2226 8134 2236 8186
rect 2260 8134 2290 8186
rect 2290 8134 2302 8186
rect 2302 8134 2316 8186
rect 2340 8134 2354 8186
rect 2354 8134 2366 8186
rect 2366 8134 2396 8186
rect 2420 8134 2430 8186
rect 2430 8134 2476 8186
rect 2180 8132 2236 8134
rect 2260 8132 2316 8134
rect 2340 8132 2396 8134
rect 2420 8132 2476 8134
rect 4628 8186 4684 8188
rect 4708 8186 4764 8188
rect 4788 8186 4844 8188
rect 4868 8186 4924 8188
rect 4628 8134 4674 8186
rect 4674 8134 4684 8186
rect 4708 8134 4738 8186
rect 4738 8134 4750 8186
rect 4750 8134 4764 8186
rect 4788 8134 4802 8186
rect 4802 8134 4814 8186
rect 4814 8134 4844 8186
rect 4868 8134 4878 8186
rect 4878 8134 4924 8186
rect 4628 8132 4684 8134
rect 4708 8132 4764 8134
rect 4788 8132 4844 8134
rect 4868 8132 4924 8134
rect 7076 8186 7132 8188
rect 7156 8186 7212 8188
rect 7236 8186 7292 8188
rect 7316 8186 7372 8188
rect 7076 8134 7122 8186
rect 7122 8134 7132 8186
rect 7156 8134 7186 8186
rect 7186 8134 7198 8186
rect 7198 8134 7212 8186
rect 7236 8134 7250 8186
rect 7250 8134 7262 8186
rect 7262 8134 7292 8186
rect 7316 8134 7326 8186
rect 7326 8134 7372 8186
rect 7076 8132 7132 8134
rect 7156 8132 7212 8134
rect 7236 8132 7292 8134
rect 7316 8132 7372 8134
rect 9524 8186 9580 8188
rect 9604 8186 9660 8188
rect 9684 8186 9740 8188
rect 9764 8186 9820 8188
rect 9524 8134 9570 8186
rect 9570 8134 9580 8186
rect 9604 8134 9634 8186
rect 9634 8134 9646 8186
rect 9646 8134 9660 8186
rect 9684 8134 9698 8186
rect 9698 8134 9710 8186
rect 9710 8134 9740 8186
rect 9764 8134 9774 8186
rect 9774 8134 9820 8186
rect 9524 8132 9580 8134
rect 9604 8132 9660 8134
rect 9684 8132 9740 8134
rect 9764 8132 9820 8134
rect 3404 7642 3460 7644
rect 3484 7642 3540 7644
rect 3564 7642 3620 7644
rect 3644 7642 3700 7644
rect 3404 7590 3450 7642
rect 3450 7590 3460 7642
rect 3484 7590 3514 7642
rect 3514 7590 3526 7642
rect 3526 7590 3540 7642
rect 3564 7590 3578 7642
rect 3578 7590 3590 7642
rect 3590 7590 3620 7642
rect 3644 7590 3654 7642
rect 3654 7590 3700 7642
rect 3404 7588 3460 7590
rect 3484 7588 3540 7590
rect 3564 7588 3620 7590
rect 3644 7588 3700 7590
rect 5852 7642 5908 7644
rect 5932 7642 5988 7644
rect 6012 7642 6068 7644
rect 6092 7642 6148 7644
rect 5852 7590 5898 7642
rect 5898 7590 5908 7642
rect 5932 7590 5962 7642
rect 5962 7590 5974 7642
rect 5974 7590 5988 7642
rect 6012 7590 6026 7642
rect 6026 7590 6038 7642
rect 6038 7590 6068 7642
rect 6092 7590 6102 7642
rect 6102 7590 6148 7642
rect 5852 7588 5908 7590
rect 5932 7588 5988 7590
rect 6012 7588 6068 7590
rect 6092 7588 6148 7590
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8540 7642 8596 7644
rect 8300 7590 8346 7642
rect 8346 7590 8356 7642
rect 8380 7590 8410 7642
rect 8410 7590 8422 7642
rect 8422 7590 8436 7642
rect 8460 7590 8474 7642
rect 8474 7590 8486 7642
rect 8486 7590 8516 7642
rect 8540 7590 8550 7642
rect 8550 7590 8596 7642
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8540 7588 8596 7590
rect 2180 7098 2236 7100
rect 2260 7098 2316 7100
rect 2340 7098 2396 7100
rect 2420 7098 2476 7100
rect 2180 7046 2226 7098
rect 2226 7046 2236 7098
rect 2260 7046 2290 7098
rect 2290 7046 2302 7098
rect 2302 7046 2316 7098
rect 2340 7046 2354 7098
rect 2354 7046 2366 7098
rect 2366 7046 2396 7098
rect 2420 7046 2430 7098
rect 2430 7046 2476 7098
rect 2180 7044 2236 7046
rect 2260 7044 2316 7046
rect 2340 7044 2396 7046
rect 2420 7044 2476 7046
rect 4628 7098 4684 7100
rect 4708 7098 4764 7100
rect 4788 7098 4844 7100
rect 4868 7098 4924 7100
rect 4628 7046 4674 7098
rect 4674 7046 4684 7098
rect 4708 7046 4738 7098
rect 4738 7046 4750 7098
rect 4750 7046 4764 7098
rect 4788 7046 4802 7098
rect 4802 7046 4814 7098
rect 4814 7046 4844 7098
rect 4868 7046 4878 7098
rect 4878 7046 4924 7098
rect 4628 7044 4684 7046
rect 4708 7044 4764 7046
rect 4788 7044 4844 7046
rect 4868 7044 4924 7046
rect 7076 7098 7132 7100
rect 7156 7098 7212 7100
rect 7236 7098 7292 7100
rect 7316 7098 7372 7100
rect 7076 7046 7122 7098
rect 7122 7046 7132 7098
rect 7156 7046 7186 7098
rect 7186 7046 7198 7098
rect 7198 7046 7212 7098
rect 7236 7046 7250 7098
rect 7250 7046 7262 7098
rect 7262 7046 7292 7098
rect 7316 7046 7326 7098
rect 7326 7046 7372 7098
rect 7076 7044 7132 7046
rect 7156 7044 7212 7046
rect 7236 7044 7292 7046
rect 7316 7044 7372 7046
rect 9524 7098 9580 7100
rect 9604 7098 9660 7100
rect 9684 7098 9740 7100
rect 9764 7098 9820 7100
rect 9524 7046 9570 7098
rect 9570 7046 9580 7098
rect 9604 7046 9634 7098
rect 9634 7046 9646 7098
rect 9646 7046 9660 7098
rect 9684 7046 9698 7098
rect 9698 7046 9710 7098
rect 9710 7046 9740 7098
rect 9764 7046 9774 7098
rect 9774 7046 9820 7098
rect 9524 7044 9580 7046
rect 9604 7044 9660 7046
rect 9684 7044 9740 7046
rect 9764 7044 9820 7046
rect 3404 6554 3460 6556
rect 3484 6554 3540 6556
rect 3564 6554 3620 6556
rect 3644 6554 3700 6556
rect 3404 6502 3450 6554
rect 3450 6502 3460 6554
rect 3484 6502 3514 6554
rect 3514 6502 3526 6554
rect 3526 6502 3540 6554
rect 3564 6502 3578 6554
rect 3578 6502 3590 6554
rect 3590 6502 3620 6554
rect 3644 6502 3654 6554
rect 3654 6502 3700 6554
rect 3404 6500 3460 6502
rect 3484 6500 3540 6502
rect 3564 6500 3620 6502
rect 3644 6500 3700 6502
rect 5852 6554 5908 6556
rect 5932 6554 5988 6556
rect 6012 6554 6068 6556
rect 6092 6554 6148 6556
rect 5852 6502 5898 6554
rect 5898 6502 5908 6554
rect 5932 6502 5962 6554
rect 5962 6502 5974 6554
rect 5974 6502 5988 6554
rect 6012 6502 6026 6554
rect 6026 6502 6038 6554
rect 6038 6502 6068 6554
rect 6092 6502 6102 6554
rect 6102 6502 6148 6554
rect 5852 6500 5908 6502
rect 5932 6500 5988 6502
rect 6012 6500 6068 6502
rect 6092 6500 6148 6502
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8540 6554 8596 6556
rect 8300 6502 8346 6554
rect 8346 6502 8356 6554
rect 8380 6502 8410 6554
rect 8410 6502 8422 6554
rect 8422 6502 8436 6554
rect 8460 6502 8474 6554
rect 8474 6502 8486 6554
rect 8486 6502 8516 6554
rect 8540 6502 8550 6554
rect 8550 6502 8596 6554
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8540 6500 8596 6502
rect 2180 6010 2236 6012
rect 2260 6010 2316 6012
rect 2340 6010 2396 6012
rect 2420 6010 2476 6012
rect 2180 5958 2226 6010
rect 2226 5958 2236 6010
rect 2260 5958 2290 6010
rect 2290 5958 2302 6010
rect 2302 5958 2316 6010
rect 2340 5958 2354 6010
rect 2354 5958 2366 6010
rect 2366 5958 2396 6010
rect 2420 5958 2430 6010
rect 2430 5958 2476 6010
rect 2180 5956 2236 5958
rect 2260 5956 2316 5958
rect 2340 5956 2396 5958
rect 2420 5956 2476 5958
rect 4628 6010 4684 6012
rect 4708 6010 4764 6012
rect 4788 6010 4844 6012
rect 4868 6010 4924 6012
rect 4628 5958 4674 6010
rect 4674 5958 4684 6010
rect 4708 5958 4738 6010
rect 4738 5958 4750 6010
rect 4750 5958 4764 6010
rect 4788 5958 4802 6010
rect 4802 5958 4814 6010
rect 4814 5958 4844 6010
rect 4868 5958 4878 6010
rect 4878 5958 4924 6010
rect 4628 5956 4684 5958
rect 4708 5956 4764 5958
rect 4788 5956 4844 5958
rect 4868 5956 4924 5958
rect 7076 6010 7132 6012
rect 7156 6010 7212 6012
rect 7236 6010 7292 6012
rect 7316 6010 7372 6012
rect 7076 5958 7122 6010
rect 7122 5958 7132 6010
rect 7156 5958 7186 6010
rect 7186 5958 7198 6010
rect 7198 5958 7212 6010
rect 7236 5958 7250 6010
rect 7250 5958 7262 6010
rect 7262 5958 7292 6010
rect 7316 5958 7326 6010
rect 7326 5958 7372 6010
rect 7076 5956 7132 5958
rect 7156 5956 7212 5958
rect 7236 5956 7292 5958
rect 7316 5956 7372 5958
rect 9524 6010 9580 6012
rect 9604 6010 9660 6012
rect 9684 6010 9740 6012
rect 9764 6010 9820 6012
rect 9524 5958 9570 6010
rect 9570 5958 9580 6010
rect 9604 5958 9634 6010
rect 9634 5958 9646 6010
rect 9646 5958 9660 6010
rect 9684 5958 9698 6010
rect 9698 5958 9710 6010
rect 9710 5958 9740 6010
rect 9764 5958 9774 6010
rect 9774 5958 9820 6010
rect 9524 5956 9580 5958
rect 9604 5956 9660 5958
rect 9684 5956 9740 5958
rect 9764 5956 9820 5958
rect 3404 5466 3460 5468
rect 3484 5466 3540 5468
rect 3564 5466 3620 5468
rect 3644 5466 3700 5468
rect 3404 5414 3450 5466
rect 3450 5414 3460 5466
rect 3484 5414 3514 5466
rect 3514 5414 3526 5466
rect 3526 5414 3540 5466
rect 3564 5414 3578 5466
rect 3578 5414 3590 5466
rect 3590 5414 3620 5466
rect 3644 5414 3654 5466
rect 3654 5414 3700 5466
rect 3404 5412 3460 5414
rect 3484 5412 3540 5414
rect 3564 5412 3620 5414
rect 3644 5412 3700 5414
rect 5852 5466 5908 5468
rect 5932 5466 5988 5468
rect 6012 5466 6068 5468
rect 6092 5466 6148 5468
rect 5852 5414 5898 5466
rect 5898 5414 5908 5466
rect 5932 5414 5962 5466
rect 5962 5414 5974 5466
rect 5974 5414 5988 5466
rect 6012 5414 6026 5466
rect 6026 5414 6038 5466
rect 6038 5414 6068 5466
rect 6092 5414 6102 5466
rect 6102 5414 6148 5466
rect 5852 5412 5908 5414
rect 5932 5412 5988 5414
rect 6012 5412 6068 5414
rect 6092 5412 6148 5414
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8540 5466 8596 5468
rect 8300 5414 8346 5466
rect 8346 5414 8356 5466
rect 8380 5414 8410 5466
rect 8410 5414 8422 5466
rect 8422 5414 8436 5466
rect 8460 5414 8474 5466
rect 8474 5414 8486 5466
rect 8486 5414 8516 5466
rect 8540 5414 8550 5466
rect 8550 5414 8596 5466
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8540 5412 8596 5414
rect 2180 4922 2236 4924
rect 2260 4922 2316 4924
rect 2340 4922 2396 4924
rect 2420 4922 2476 4924
rect 2180 4870 2226 4922
rect 2226 4870 2236 4922
rect 2260 4870 2290 4922
rect 2290 4870 2302 4922
rect 2302 4870 2316 4922
rect 2340 4870 2354 4922
rect 2354 4870 2366 4922
rect 2366 4870 2396 4922
rect 2420 4870 2430 4922
rect 2430 4870 2476 4922
rect 2180 4868 2236 4870
rect 2260 4868 2316 4870
rect 2340 4868 2396 4870
rect 2420 4868 2476 4870
rect 4628 4922 4684 4924
rect 4708 4922 4764 4924
rect 4788 4922 4844 4924
rect 4868 4922 4924 4924
rect 4628 4870 4674 4922
rect 4674 4870 4684 4922
rect 4708 4870 4738 4922
rect 4738 4870 4750 4922
rect 4750 4870 4764 4922
rect 4788 4870 4802 4922
rect 4802 4870 4814 4922
rect 4814 4870 4844 4922
rect 4868 4870 4878 4922
rect 4878 4870 4924 4922
rect 4628 4868 4684 4870
rect 4708 4868 4764 4870
rect 4788 4868 4844 4870
rect 4868 4868 4924 4870
rect 7076 4922 7132 4924
rect 7156 4922 7212 4924
rect 7236 4922 7292 4924
rect 7316 4922 7372 4924
rect 7076 4870 7122 4922
rect 7122 4870 7132 4922
rect 7156 4870 7186 4922
rect 7186 4870 7198 4922
rect 7198 4870 7212 4922
rect 7236 4870 7250 4922
rect 7250 4870 7262 4922
rect 7262 4870 7292 4922
rect 7316 4870 7326 4922
rect 7326 4870 7372 4922
rect 7076 4868 7132 4870
rect 7156 4868 7212 4870
rect 7236 4868 7292 4870
rect 7316 4868 7372 4870
rect 9524 4922 9580 4924
rect 9604 4922 9660 4924
rect 9684 4922 9740 4924
rect 9764 4922 9820 4924
rect 9524 4870 9570 4922
rect 9570 4870 9580 4922
rect 9604 4870 9634 4922
rect 9634 4870 9646 4922
rect 9646 4870 9660 4922
rect 9684 4870 9698 4922
rect 9698 4870 9710 4922
rect 9710 4870 9740 4922
rect 9764 4870 9774 4922
rect 9774 4870 9820 4922
rect 9524 4868 9580 4870
rect 9604 4868 9660 4870
rect 9684 4868 9740 4870
rect 9764 4868 9820 4870
rect 3404 4378 3460 4380
rect 3484 4378 3540 4380
rect 3564 4378 3620 4380
rect 3644 4378 3700 4380
rect 3404 4326 3450 4378
rect 3450 4326 3460 4378
rect 3484 4326 3514 4378
rect 3514 4326 3526 4378
rect 3526 4326 3540 4378
rect 3564 4326 3578 4378
rect 3578 4326 3590 4378
rect 3590 4326 3620 4378
rect 3644 4326 3654 4378
rect 3654 4326 3700 4378
rect 3404 4324 3460 4326
rect 3484 4324 3540 4326
rect 3564 4324 3620 4326
rect 3644 4324 3700 4326
rect 2180 3834 2236 3836
rect 2260 3834 2316 3836
rect 2340 3834 2396 3836
rect 2420 3834 2476 3836
rect 2180 3782 2226 3834
rect 2226 3782 2236 3834
rect 2260 3782 2290 3834
rect 2290 3782 2302 3834
rect 2302 3782 2316 3834
rect 2340 3782 2354 3834
rect 2354 3782 2366 3834
rect 2366 3782 2396 3834
rect 2420 3782 2430 3834
rect 2430 3782 2476 3834
rect 2180 3780 2236 3782
rect 2260 3780 2316 3782
rect 2340 3780 2396 3782
rect 2420 3780 2476 3782
rect 2180 2746 2236 2748
rect 2260 2746 2316 2748
rect 2340 2746 2396 2748
rect 2420 2746 2476 2748
rect 2180 2694 2226 2746
rect 2226 2694 2236 2746
rect 2260 2694 2290 2746
rect 2290 2694 2302 2746
rect 2302 2694 2316 2746
rect 2340 2694 2354 2746
rect 2354 2694 2366 2746
rect 2366 2694 2396 2746
rect 2420 2694 2430 2746
rect 2430 2694 2476 2746
rect 2180 2692 2236 2694
rect 2260 2692 2316 2694
rect 2340 2692 2396 2694
rect 2420 2692 2476 2694
rect 3404 3290 3460 3292
rect 3484 3290 3540 3292
rect 3564 3290 3620 3292
rect 3644 3290 3700 3292
rect 3404 3238 3450 3290
rect 3450 3238 3460 3290
rect 3484 3238 3514 3290
rect 3514 3238 3526 3290
rect 3526 3238 3540 3290
rect 3564 3238 3578 3290
rect 3578 3238 3590 3290
rect 3590 3238 3620 3290
rect 3644 3238 3654 3290
rect 3654 3238 3700 3290
rect 3404 3236 3460 3238
rect 3484 3236 3540 3238
rect 3564 3236 3620 3238
rect 3644 3236 3700 3238
rect 3404 2202 3460 2204
rect 3484 2202 3540 2204
rect 3564 2202 3620 2204
rect 3644 2202 3700 2204
rect 3404 2150 3450 2202
rect 3450 2150 3460 2202
rect 3484 2150 3514 2202
rect 3514 2150 3526 2202
rect 3526 2150 3540 2202
rect 3564 2150 3578 2202
rect 3578 2150 3590 2202
rect 3590 2150 3620 2202
rect 3644 2150 3654 2202
rect 3654 2150 3700 2202
rect 3404 2148 3460 2150
rect 3484 2148 3540 2150
rect 3564 2148 3620 2150
rect 3644 2148 3700 2150
rect 5852 4378 5908 4380
rect 5932 4378 5988 4380
rect 6012 4378 6068 4380
rect 6092 4378 6148 4380
rect 5852 4326 5898 4378
rect 5898 4326 5908 4378
rect 5932 4326 5962 4378
rect 5962 4326 5974 4378
rect 5974 4326 5988 4378
rect 6012 4326 6026 4378
rect 6026 4326 6038 4378
rect 6038 4326 6068 4378
rect 6092 4326 6102 4378
rect 6102 4326 6148 4378
rect 5852 4324 5908 4326
rect 5932 4324 5988 4326
rect 6012 4324 6068 4326
rect 6092 4324 6148 4326
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8540 4378 8596 4380
rect 8300 4326 8346 4378
rect 8346 4326 8356 4378
rect 8380 4326 8410 4378
rect 8410 4326 8422 4378
rect 8422 4326 8436 4378
rect 8460 4326 8474 4378
rect 8474 4326 8486 4378
rect 8486 4326 8516 4378
rect 8540 4326 8550 4378
rect 8550 4326 8596 4378
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8540 4324 8596 4326
rect 4628 3834 4684 3836
rect 4708 3834 4764 3836
rect 4788 3834 4844 3836
rect 4868 3834 4924 3836
rect 4628 3782 4674 3834
rect 4674 3782 4684 3834
rect 4708 3782 4738 3834
rect 4738 3782 4750 3834
rect 4750 3782 4764 3834
rect 4788 3782 4802 3834
rect 4802 3782 4814 3834
rect 4814 3782 4844 3834
rect 4868 3782 4878 3834
rect 4878 3782 4924 3834
rect 4628 3780 4684 3782
rect 4708 3780 4764 3782
rect 4788 3780 4844 3782
rect 4868 3780 4924 3782
rect 4628 2746 4684 2748
rect 4708 2746 4764 2748
rect 4788 2746 4844 2748
rect 4868 2746 4924 2748
rect 4628 2694 4674 2746
rect 4674 2694 4684 2746
rect 4708 2694 4738 2746
rect 4738 2694 4750 2746
rect 4750 2694 4764 2746
rect 4788 2694 4802 2746
rect 4802 2694 4814 2746
rect 4814 2694 4844 2746
rect 4868 2694 4878 2746
rect 4878 2694 4924 2746
rect 4628 2692 4684 2694
rect 4708 2692 4764 2694
rect 4788 2692 4844 2694
rect 4868 2692 4924 2694
rect 5852 3290 5908 3292
rect 5932 3290 5988 3292
rect 6012 3290 6068 3292
rect 6092 3290 6148 3292
rect 5852 3238 5898 3290
rect 5898 3238 5908 3290
rect 5932 3238 5962 3290
rect 5962 3238 5974 3290
rect 5974 3238 5988 3290
rect 6012 3238 6026 3290
rect 6026 3238 6038 3290
rect 6038 3238 6068 3290
rect 6092 3238 6102 3290
rect 6102 3238 6148 3290
rect 5852 3236 5908 3238
rect 5932 3236 5988 3238
rect 6012 3236 6068 3238
rect 6092 3236 6148 3238
rect 5852 2202 5908 2204
rect 5932 2202 5988 2204
rect 6012 2202 6068 2204
rect 6092 2202 6148 2204
rect 5852 2150 5898 2202
rect 5898 2150 5908 2202
rect 5932 2150 5962 2202
rect 5962 2150 5974 2202
rect 5974 2150 5988 2202
rect 6012 2150 6026 2202
rect 6026 2150 6038 2202
rect 6038 2150 6068 2202
rect 6092 2150 6102 2202
rect 6102 2150 6148 2202
rect 5852 2148 5908 2150
rect 5932 2148 5988 2150
rect 6012 2148 6068 2150
rect 6092 2148 6148 2150
rect 7076 3834 7132 3836
rect 7156 3834 7212 3836
rect 7236 3834 7292 3836
rect 7316 3834 7372 3836
rect 7076 3782 7122 3834
rect 7122 3782 7132 3834
rect 7156 3782 7186 3834
rect 7186 3782 7198 3834
rect 7198 3782 7212 3834
rect 7236 3782 7250 3834
rect 7250 3782 7262 3834
rect 7262 3782 7292 3834
rect 7316 3782 7326 3834
rect 7326 3782 7372 3834
rect 7076 3780 7132 3782
rect 7156 3780 7212 3782
rect 7236 3780 7292 3782
rect 7316 3780 7372 3782
rect 7076 2746 7132 2748
rect 7156 2746 7212 2748
rect 7236 2746 7292 2748
rect 7316 2746 7372 2748
rect 7076 2694 7122 2746
rect 7122 2694 7132 2746
rect 7156 2694 7186 2746
rect 7186 2694 7198 2746
rect 7198 2694 7212 2746
rect 7236 2694 7250 2746
rect 7250 2694 7262 2746
rect 7262 2694 7292 2746
rect 7316 2694 7326 2746
rect 7326 2694 7372 2746
rect 7076 2692 7132 2694
rect 7156 2692 7212 2694
rect 7236 2692 7292 2694
rect 7316 2692 7372 2694
rect 9524 3834 9580 3836
rect 9604 3834 9660 3836
rect 9684 3834 9740 3836
rect 9764 3834 9820 3836
rect 9524 3782 9570 3834
rect 9570 3782 9580 3834
rect 9604 3782 9634 3834
rect 9634 3782 9646 3834
rect 9646 3782 9660 3834
rect 9684 3782 9698 3834
rect 9698 3782 9710 3834
rect 9710 3782 9740 3834
rect 9764 3782 9774 3834
rect 9774 3782 9820 3834
rect 9524 3780 9580 3782
rect 9604 3780 9660 3782
rect 9684 3780 9740 3782
rect 9764 3780 9820 3782
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8540 3290 8596 3292
rect 8300 3238 8346 3290
rect 8346 3238 8356 3290
rect 8380 3238 8410 3290
rect 8410 3238 8422 3290
rect 8422 3238 8436 3290
rect 8460 3238 8474 3290
rect 8474 3238 8486 3290
rect 8486 3238 8516 3290
rect 8540 3238 8550 3290
rect 8550 3238 8596 3290
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8540 3236 8596 3238
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8540 2202 8596 2204
rect 8300 2150 8346 2202
rect 8346 2150 8356 2202
rect 8380 2150 8410 2202
rect 8410 2150 8422 2202
rect 8422 2150 8436 2202
rect 8460 2150 8474 2202
rect 8474 2150 8486 2202
rect 8486 2150 8516 2202
rect 8540 2150 8550 2202
rect 8550 2150 8596 2202
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8540 2148 8596 2150
rect 9524 2746 9580 2748
rect 9604 2746 9660 2748
rect 9684 2746 9740 2748
rect 9764 2746 9820 2748
rect 9524 2694 9570 2746
rect 9570 2694 9580 2746
rect 9604 2694 9634 2746
rect 9634 2694 9646 2746
rect 9646 2694 9660 2746
rect 9684 2694 9698 2746
rect 9698 2694 9710 2746
rect 9710 2694 9740 2746
rect 9764 2694 9774 2746
rect 9774 2694 9820 2746
rect 9524 2692 9580 2694
rect 9604 2692 9660 2694
rect 9684 2692 9740 2694
rect 9764 2692 9820 2694
<< metal3 >>
rect 2170 11456 2486 11457
rect 2170 11392 2176 11456
rect 2240 11392 2256 11456
rect 2320 11392 2336 11456
rect 2400 11392 2416 11456
rect 2480 11392 2486 11456
rect 2170 11391 2486 11392
rect 4618 11456 4934 11457
rect 4618 11392 4624 11456
rect 4688 11392 4704 11456
rect 4768 11392 4784 11456
rect 4848 11392 4864 11456
rect 4928 11392 4934 11456
rect 4618 11391 4934 11392
rect 7066 11456 7382 11457
rect 7066 11392 7072 11456
rect 7136 11392 7152 11456
rect 7216 11392 7232 11456
rect 7296 11392 7312 11456
rect 7376 11392 7382 11456
rect 7066 11391 7382 11392
rect 9514 11456 9830 11457
rect 9514 11392 9520 11456
rect 9584 11392 9600 11456
rect 9664 11392 9680 11456
rect 9744 11392 9760 11456
rect 9824 11392 9830 11456
rect 9514 11391 9830 11392
rect 3394 10912 3710 10913
rect 3394 10848 3400 10912
rect 3464 10848 3480 10912
rect 3544 10848 3560 10912
rect 3624 10848 3640 10912
rect 3704 10848 3710 10912
rect 3394 10847 3710 10848
rect 5842 10912 6158 10913
rect 5842 10848 5848 10912
rect 5912 10848 5928 10912
rect 5992 10848 6008 10912
rect 6072 10848 6088 10912
rect 6152 10848 6158 10912
rect 5842 10847 6158 10848
rect 8290 10912 8606 10913
rect 8290 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8536 10912
rect 8600 10848 8606 10912
rect 8290 10847 8606 10848
rect 2170 10368 2486 10369
rect 2170 10304 2176 10368
rect 2240 10304 2256 10368
rect 2320 10304 2336 10368
rect 2400 10304 2416 10368
rect 2480 10304 2486 10368
rect 2170 10303 2486 10304
rect 4618 10368 4934 10369
rect 4618 10304 4624 10368
rect 4688 10304 4704 10368
rect 4768 10304 4784 10368
rect 4848 10304 4864 10368
rect 4928 10304 4934 10368
rect 4618 10303 4934 10304
rect 7066 10368 7382 10369
rect 7066 10304 7072 10368
rect 7136 10304 7152 10368
rect 7216 10304 7232 10368
rect 7296 10304 7312 10368
rect 7376 10304 7382 10368
rect 7066 10303 7382 10304
rect 9514 10368 9830 10369
rect 9514 10304 9520 10368
rect 9584 10304 9600 10368
rect 9664 10304 9680 10368
rect 9744 10304 9760 10368
rect 9824 10304 9830 10368
rect 9514 10303 9830 10304
rect 3394 9824 3710 9825
rect 3394 9760 3400 9824
rect 3464 9760 3480 9824
rect 3544 9760 3560 9824
rect 3624 9760 3640 9824
rect 3704 9760 3710 9824
rect 3394 9759 3710 9760
rect 5842 9824 6158 9825
rect 5842 9760 5848 9824
rect 5912 9760 5928 9824
rect 5992 9760 6008 9824
rect 6072 9760 6088 9824
rect 6152 9760 6158 9824
rect 5842 9759 6158 9760
rect 8290 9824 8606 9825
rect 8290 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8536 9824
rect 8600 9760 8606 9824
rect 8290 9759 8606 9760
rect 2170 9280 2486 9281
rect 2170 9216 2176 9280
rect 2240 9216 2256 9280
rect 2320 9216 2336 9280
rect 2400 9216 2416 9280
rect 2480 9216 2486 9280
rect 2170 9215 2486 9216
rect 4618 9280 4934 9281
rect 4618 9216 4624 9280
rect 4688 9216 4704 9280
rect 4768 9216 4784 9280
rect 4848 9216 4864 9280
rect 4928 9216 4934 9280
rect 4618 9215 4934 9216
rect 7066 9280 7382 9281
rect 7066 9216 7072 9280
rect 7136 9216 7152 9280
rect 7216 9216 7232 9280
rect 7296 9216 7312 9280
rect 7376 9216 7382 9280
rect 7066 9215 7382 9216
rect 9514 9280 9830 9281
rect 9514 9216 9520 9280
rect 9584 9216 9600 9280
rect 9664 9216 9680 9280
rect 9744 9216 9760 9280
rect 9824 9216 9830 9280
rect 9514 9215 9830 9216
rect 3394 8736 3710 8737
rect 3394 8672 3400 8736
rect 3464 8672 3480 8736
rect 3544 8672 3560 8736
rect 3624 8672 3640 8736
rect 3704 8672 3710 8736
rect 3394 8671 3710 8672
rect 5842 8736 6158 8737
rect 5842 8672 5848 8736
rect 5912 8672 5928 8736
rect 5992 8672 6008 8736
rect 6072 8672 6088 8736
rect 6152 8672 6158 8736
rect 5842 8671 6158 8672
rect 8290 8736 8606 8737
rect 8290 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8536 8736
rect 8600 8672 8606 8736
rect 8290 8671 8606 8672
rect 2170 8192 2486 8193
rect 2170 8128 2176 8192
rect 2240 8128 2256 8192
rect 2320 8128 2336 8192
rect 2400 8128 2416 8192
rect 2480 8128 2486 8192
rect 2170 8127 2486 8128
rect 4618 8192 4934 8193
rect 4618 8128 4624 8192
rect 4688 8128 4704 8192
rect 4768 8128 4784 8192
rect 4848 8128 4864 8192
rect 4928 8128 4934 8192
rect 4618 8127 4934 8128
rect 7066 8192 7382 8193
rect 7066 8128 7072 8192
rect 7136 8128 7152 8192
rect 7216 8128 7232 8192
rect 7296 8128 7312 8192
rect 7376 8128 7382 8192
rect 7066 8127 7382 8128
rect 9514 8192 9830 8193
rect 9514 8128 9520 8192
rect 9584 8128 9600 8192
rect 9664 8128 9680 8192
rect 9744 8128 9760 8192
rect 9824 8128 9830 8192
rect 9514 8127 9830 8128
rect 3394 7648 3710 7649
rect 3394 7584 3400 7648
rect 3464 7584 3480 7648
rect 3544 7584 3560 7648
rect 3624 7584 3640 7648
rect 3704 7584 3710 7648
rect 3394 7583 3710 7584
rect 5842 7648 6158 7649
rect 5842 7584 5848 7648
rect 5912 7584 5928 7648
rect 5992 7584 6008 7648
rect 6072 7584 6088 7648
rect 6152 7584 6158 7648
rect 5842 7583 6158 7584
rect 8290 7648 8606 7649
rect 8290 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8536 7648
rect 8600 7584 8606 7648
rect 8290 7583 8606 7584
rect 2170 7104 2486 7105
rect 2170 7040 2176 7104
rect 2240 7040 2256 7104
rect 2320 7040 2336 7104
rect 2400 7040 2416 7104
rect 2480 7040 2486 7104
rect 2170 7039 2486 7040
rect 4618 7104 4934 7105
rect 4618 7040 4624 7104
rect 4688 7040 4704 7104
rect 4768 7040 4784 7104
rect 4848 7040 4864 7104
rect 4928 7040 4934 7104
rect 4618 7039 4934 7040
rect 7066 7104 7382 7105
rect 7066 7040 7072 7104
rect 7136 7040 7152 7104
rect 7216 7040 7232 7104
rect 7296 7040 7312 7104
rect 7376 7040 7382 7104
rect 7066 7039 7382 7040
rect 9514 7104 9830 7105
rect 9514 7040 9520 7104
rect 9584 7040 9600 7104
rect 9664 7040 9680 7104
rect 9744 7040 9760 7104
rect 9824 7040 9830 7104
rect 9514 7039 9830 7040
rect 3394 6560 3710 6561
rect 3394 6496 3400 6560
rect 3464 6496 3480 6560
rect 3544 6496 3560 6560
rect 3624 6496 3640 6560
rect 3704 6496 3710 6560
rect 3394 6495 3710 6496
rect 5842 6560 6158 6561
rect 5842 6496 5848 6560
rect 5912 6496 5928 6560
rect 5992 6496 6008 6560
rect 6072 6496 6088 6560
rect 6152 6496 6158 6560
rect 5842 6495 6158 6496
rect 8290 6560 8606 6561
rect 8290 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8536 6560
rect 8600 6496 8606 6560
rect 8290 6495 8606 6496
rect 2170 6016 2486 6017
rect 2170 5952 2176 6016
rect 2240 5952 2256 6016
rect 2320 5952 2336 6016
rect 2400 5952 2416 6016
rect 2480 5952 2486 6016
rect 2170 5951 2486 5952
rect 4618 6016 4934 6017
rect 4618 5952 4624 6016
rect 4688 5952 4704 6016
rect 4768 5952 4784 6016
rect 4848 5952 4864 6016
rect 4928 5952 4934 6016
rect 4618 5951 4934 5952
rect 7066 6016 7382 6017
rect 7066 5952 7072 6016
rect 7136 5952 7152 6016
rect 7216 5952 7232 6016
rect 7296 5952 7312 6016
rect 7376 5952 7382 6016
rect 7066 5951 7382 5952
rect 9514 6016 9830 6017
rect 9514 5952 9520 6016
rect 9584 5952 9600 6016
rect 9664 5952 9680 6016
rect 9744 5952 9760 6016
rect 9824 5952 9830 6016
rect 9514 5951 9830 5952
rect 3394 5472 3710 5473
rect 3394 5408 3400 5472
rect 3464 5408 3480 5472
rect 3544 5408 3560 5472
rect 3624 5408 3640 5472
rect 3704 5408 3710 5472
rect 3394 5407 3710 5408
rect 5842 5472 6158 5473
rect 5842 5408 5848 5472
rect 5912 5408 5928 5472
rect 5992 5408 6008 5472
rect 6072 5408 6088 5472
rect 6152 5408 6158 5472
rect 5842 5407 6158 5408
rect 8290 5472 8606 5473
rect 8290 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8536 5472
rect 8600 5408 8606 5472
rect 8290 5407 8606 5408
rect 2170 4928 2486 4929
rect 2170 4864 2176 4928
rect 2240 4864 2256 4928
rect 2320 4864 2336 4928
rect 2400 4864 2416 4928
rect 2480 4864 2486 4928
rect 2170 4863 2486 4864
rect 4618 4928 4934 4929
rect 4618 4864 4624 4928
rect 4688 4864 4704 4928
rect 4768 4864 4784 4928
rect 4848 4864 4864 4928
rect 4928 4864 4934 4928
rect 4618 4863 4934 4864
rect 7066 4928 7382 4929
rect 7066 4864 7072 4928
rect 7136 4864 7152 4928
rect 7216 4864 7232 4928
rect 7296 4864 7312 4928
rect 7376 4864 7382 4928
rect 7066 4863 7382 4864
rect 9514 4928 9830 4929
rect 9514 4864 9520 4928
rect 9584 4864 9600 4928
rect 9664 4864 9680 4928
rect 9744 4864 9760 4928
rect 9824 4864 9830 4928
rect 9514 4863 9830 4864
rect 3394 4384 3710 4385
rect 3394 4320 3400 4384
rect 3464 4320 3480 4384
rect 3544 4320 3560 4384
rect 3624 4320 3640 4384
rect 3704 4320 3710 4384
rect 3394 4319 3710 4320
rect 5842 4384 6158 4385
rect 5842 4320 5848 4384
rect 5912 4320 5928 4384
rect 5992 4320 6008 4384
rect 6072 4320 6088 4384
rect 6152 4320 6158 4384
rect 5842 4319 6158 4320
rect 8290 4384 8606 4385
rect 8290 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8536 4384
rect 8600 4320 8606 4384
rect 8290 4319 8606 4320
rect 2170 3840 2486 3841
rect 2170 3776 2176 3840
rect 2240 3776 2256 3840
rect 2320 3776 2336 3840
rect 2400 3776 2416 3840
rect 2480 3776 2486 3840
rect 2170 3775 2486 3776
rect 4618 3840 4934 3841
rect 4618 3776 4624 3840
rect 4688 3776 4704 3840
rect 4768 3776 4784 3840
rect 4848 3776 4864 3840
rect 4928 3776 4934 3840
rect 4618 3775 4934 3776
rect 7066 3840 7382 3841
rect 7066 3776 7072 3840
rect 7136 3776 7152 3840
rect 7216 3776 7232 3840
rect 7296 3776 7312 3840
rect 7376 3776 7382 3840
rect 7066 3775 7382 3776
rect 9514 3840 9830 3841
rect 9514 3776 9520 3840
rect 9584 3776 9600 3840
rect 9664 3776 9680 3840
rect 9744 3776 9760 3840
rect 9824 3776 9830 3840
rect 9514 3775 9830 3776
rect 3394 3296 3710 3297
rect 3394 3232 3400 3296
rect 3464 3232 3480 3296
rect 3544 3232 3560 3296
rect 3624 3232 3640 3296
rect 3704 3232 3710 3296
rect 3394 3231 3710 3232
rect 5842 3296 6158 3297
rect 5842 3232 5848 3296
rect 5912 3232 5928 3296
rect 5992 3232 6008 3296
rect 6072 3232 6088 3296
rect 6152 3232 6158 3296
rect 5842 3231 6158 3232
rect 8290 3296 8606 3297
rect 8290 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8536 3296
rect 8600 3232 8606 3296
rect 8290 3231 8606 3232
rect 2170 2752 2486 2753
rect 2170 2688 2176 2752
rect 2240 2688 2256 2752
rect 2320 2688 2336 2752
rect 2400 2688 2416 2752
rect 2480 2688 2486 2752
rect 2170 2687 2486 2688
rect 4618 2752 4934 2753
rect 4618 2688 4624 2752
rect 4688 2688 4704 2752
rect 4768 2688 4784 2752
rect 4848 2688 4864 2752
rect 4928 2688 4934 2752
rect 4618 2687 4934 2688
rect 7066 2752 7382 2753
rect 7066 2688 7072 2752
rect 7136 2688 7152 2752
rect 7216 2688 7232 2752
rect 7296 2688 7312 2752
rect 7376 2688 7382 2752
rect 7066 2687 7382 2688
rect 9514 2752 9830 2753
rect 9514 2688 9520 2752
rect 9584 2688 9600 2752
rect 9664 2688 9680 2752
rect 9744 2688 9760 2752
rect 9824 2688 9830 2752
rect 9514 2687 9830 2688
rect 3394 2208 3710 2209
rect 3394 2144 3400 2208
rect 3464 2144 3480 2208
rect 3544 2144 3560 2208
rect 3624 2144 3640 2208
rect 3704 2144 3710 2208
rect 3394 2143 3710 2144
rect 5842 2208 6158 2209
rect 5842 2144 5848 2208
rect 5912 2144 5928 2208
rect 5992 2144 6008 2208
rect 6072 2144 6088 2208
rect 6152 2144 6158 2208
rect 5842 2143 6158 2144
rect 8290 2208 8606 2209
rect 8290 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8536 2208
rect 8600 2144 8606 2208
rect 8290 2143 8606 2144
<< via3 >>
rect 2176 11452 2240 11456
rect 2176 11396 2180 11452
rect 2180 11396 2236 11452
rect 2236 11396 2240 11452
rect 2176 11392 2240 11396
rect 2256 11452 2320 11456
rect 2256 11396 2260 11452
rect 2260 11396 2316 11452
rect 2316 11396 2320 11452
rect 2256 11392 2320 11396
rect 2336 11452 2400 11456
rect 2336 11396 2340 11452
rect 2340 11396 2396 11452
rect 2396 11396 2400 11452
rect 2336 11392 2400 11396
rect 2416 11452 2480 11456
rect 2416 11396 2420 11452
rect 2420 11396 2476 11452
rect 2476 11396 2480 11452
rect 2416 11392 2480 11396
rect 4624 11452 4688 11456
rect 4624 11396 4628 11452
rect 4628 11396 4684 11452
rect 4684 11396 4688 11452
rect 4624 11392 4688 11396
rect 4704 11452 4768 11456
rect 4704 11396 4708 11452
rect 4708 11396 4764 11452
rect 4764 11396 4768 11452
rect 4704 11392 4768 11396
rect 4784 11452 4848 11456
rect 4784 11396 4788 11452
rect 4788 11396 4844 11452
rect 4844 11396 4848 11452
rect 4784 11392 4848 11396
rect 4864 11452 4928 11456
rect 4864 11396 4868 11452
rect 4868 11396 4924 11452
rect 4924 11396 4928 11452
rect 4864 11392 4928 11396
rect 7072 11452 7136 11456
rect 7072 11396 7076 11452
rect 7076 11396 7132 11452
rect 7132 11396 7136 11452
rect 7072 11392 7136 11396
rect 7152 11452 7216 11456
rect 7152 11396 7156 11452
rect 7156 11396 7212 11452
rect 7212 11396 7216 11452
rect 7152 11392 7216 11396
rect 7232 11452 7296 11456
rect 7232 11396 7236 11452
rect 7236 11396 7292 11452
rect 7292 11396 7296 11452
rect 7232 11392 7296 11396
rect 7312 11452 7376 11456
rect 7312 11396 7316 11452
rect 7316 11396 7372 11452
rect 7372 11396 7376 11452
rect 7312 11392 7376 11396
rect 9520 11452 9584 11456
rect 9520 11396 9524 11452
rect 9524 11396 9580 11452
rect 9580 11396 9584 11452
rect 9520 11392 9584 11396
rect 9600 11452 9664 11456
rect 9600 11396 9604 11452
rect 9604 11396 9660 11452
rect 9660 11396 9664 11452
rect 9600 11392 9664 11396
rect 9680 11452 9744 11456
rect 9680 11396 9684 11452
rect 9684 11396 9740 11452
rect 9740 11396 9744 11452
rect 9680 11392 9744 11396
rect 9760 11452 9824 11456
rect 9760 11396 9764 11452
rect 9764 11396 9820 11452
rect 9820 11396 9824 11452
rect 9760 11392 9824 11396
rect 3400 10908 3464 10912
rect 3400 10852 3404 10908
rect 3404 10852 3460 10908
rect 3460 10852 3464 10908
rect 3400 10848 3464 10852
rect 3480 10908 3544 10912
rect 3480 10852 3484 10908
rect 3484 10852 3540 10908
rect 3540 10852 3544 10908
rect 3480 10848 3544 10852
rect 3560 10908 3624 10912
rect 3560 10852 3564 10908
rect 3564 10852 3620 10908
rect 3620 10852 3624 10908
rect 3560 10848 3624 10852
rect 3640 10908 3704 10912
rect 3640 10852 3644 10908
rect 3644 10852 3700 10908
rect 3700 10852 3704 10908
rect 3640 10848 3704 10852
rect 5848 10908 5912 10912
rect 5848 10852 5852 10908
rect 5852 10852 5908 10908
rect 5908 10852 5912 10908
rect 5848 10848 5912 10852
rect 5928 10908 5992 10912
rect 5928 10852 5932 10908
rect 5932 10852 5988 10908
rect 5988 10852 5992 10908
rect 5928 10848 5992 10852
rect 6008 10908 6072 10912
rect 6008 10852 6012 10908
rect 6012 10852 6068 10908
rect 6068 10852 6072 10908
rect 6008 10848 6072 10852
rect 6088 10908 6152 10912
rect 6088 10852 6092 10908
rect 6092 10852 6148 10908
rect 6148 10852 6152 10908
rect 6088 10848 6152 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 8536 10908 8600 10912
rect 8536 10852 8540 10908
rect 8540 10852 8596 10908
rect 8596 10852 8600 10908
rect 8536 10848 8600 10852
rect 2176 10364 2240 10368
rect 2176 10308 2180 10364
rect 2180 10308 2236 10364
rect 2236 10308 2240 10364
rect 2176 10304 2240 10308
rect 2256 10364 2320 10368
rect 2256 10308 2260 10364
rect 2260 10308 2316 10364
rect 2316 10308 2320 10364
rect 2256 10304 2320 10308
rect 2336 10364 2400 10368
rect 2336 10308 2340 10364
rect 2340 10308 2396 10364
rect 2396 10308 2400 10364
rect 2336 10304 2400 10308
rect 2416 10364 2480 10368
rect 2416 10308 2420 10364
rect 2420 10308 2476 10364
rect 2476 10308 2480 10364
rect 2416 10304 2480 10308
rect 4624 10364 4688 10368
rect 4624 10308 4628 10364
rect 4628 10308 4684 10364
rect 4684 10308 4688 10364
rect 4624 10304 4688 10308
rect 4704 10364 4768 10368
rect 4704 10308 4708 10364
rect 4708 10308 4764 10364
rect 4764 10308 4768 10364
rect 4704 10304 4768 10308
rect 4784 10364 4848 10368
rect 4784 10308 4788 10364
rect 4788 10308 4844 10364
rect 4844 10308 4848 10364
rect 4784 10304 4848 10308
rect 4864 10364 4928 10368
rect 4864 10308 4868 10364
rect 4868 10308 4924 10364
rect 4924 10308 4928 10364
rect 4864 10304 4928 10308
rect 7072 10364 7136 10368
rect 7072 10308 7076 10364
rect 7076 10308 7132 10364
rect 7132 10308 7136 10364
rect 7072 10304 7136 10308
rect 7152 10364 7216 10368
rect 7152 10308 7156 10364
rect 7156 10308 7212 10364
rect 7212 10308 7216 10364
rect 7152 10304 7216 10308
rect 7232 10364 7296 10368
rect 7232 10308 7236 10364
rect 7236 10308 7292 10364
rect 7292 10308 7296 10364
rect 7232 10304 7296 10308
rect 7312 10364 7376 10368
rect 7312 10308 7316 10364
rect 7316 10308 7372 10364
rect 7372 10308 7376 10364
rect 7312 10304 7376 10308
rect 9520 10364 9584 10368
rect 9520 10308 9524 10364
rect 9524 10308 9580 10364
rect 9580 10308 9584 10364
rect 9520 10304 9584 10308
rect 9600 10364 9664 10368
rect 9600 10308 9604 10364
rect 9604 10308 9660 10364
rect 9660 10308 9664 10364
rect 9600 10304 9664 10308
rect 9680 10364 9744 10368
rect 9680 10308 9684 10364
rect 9684 10308 9740 10364
rect 9740 10308 9744 10364
rect 9680 10304 9744 10308
rect 9760 10364 9824 10368
rect 9760 10308 9764 10364
rect 9764 10308 9820 10364
rect 9820 10308 9824 10364
rect 9760 10304 9824 10308
rect 3400 9820 3464 9824
rect 3400 9764 3404 9820
rect 3404 9764 3460 9820
rect 3460 9764 3464 9820
rect 3400 9760 3464 9764
rect 3480 9820 3544 9824
rect 3480 9764 3484 9820
rect 3484 9764 3540 9820
rect 3540 9764 3544 9820
rect 3480 9760 3544 9764
rect 3560 9820 3624 9824
rect 3560 9764 3564 9820
rect 3564 9764 3620 9820
rect 3620 9764 3624 9820
rect 3560 9760 3624 9764
rect 3640 9820 3704 9824
rect 3640 9764 3644 9820
rect 3644 9764 3700 9820
rect 3700 9764 3704 9820
rect 3640 9760 3704 9764
rect 5848 9820 5912 9824
rect 5848 9764 5852 9820
rect 5852 9764 5908 9820
rect 5908 9764 5912 9820
rect 5848 9760 5912 9764
rect 5928 9820 5992 9824
rect 5928 9764 5932 9820
rect 5932 9764 5988 9820
rect 5988 9764 5992 9820
rect 5928 9760 5992 9764
rect 6008 9820 6072 9824
rect 6008 9764 6012 9820
rect 6012 9764 6068 9820
rect 6068 9764 6072 9820
rect 6008 9760 6072 9764
rect 6088 9820 6152 9824
rect 6088 9764 6092 9820
rect 6092 9764 6148 9820
rect 6148 9764 6152 9820
rect 6088 9760 6152 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 8536 9820 8600 9824
rect 8536 9764 8540 9820
rect 8540 9764 8596 9820
rect 8596 9764 8600 9820
rect 8536 9760 8600 9764
rect 2176 9276 2240 9280
rect 2176 9220 2180 9276
rect 2180 9220 2236 9276
rect 2236 9220 2240 9276
rect 2176 9216 2240 9220
rect 2256 9276 2320 9280
rect 2256 9220 2260 9276
rect 2260 9220 2316 9276
rect 2316 9220 2320 9276
rect 2256 9216 2320 9220
rect 2336 9276 2400 9280
rect 2336 9220 2340 9276
rect 2340 9220 2396 9276
rect 2396 9220 2400 9276
rect 2336 9216 2400 9220
rect 2416 9276 2480 9280
rect 2416 9220 2420 9276
rect 2420 9220 2476 9276
rect 2476 9220 2480 9276
rect 2416 9216 2480 9220
rect 4624 9276 4688 9280
rect 4624 9220 4628 9276
rect 4628 9220 4684 9276
rect 4684 9220 4688 9276
rect 4624 9216 4688 9220
rect 4704 9276 4768 9280
rect 4704 9220 4708 9276
rect 4708 9220 4764 9276
rect 4764 9220 4768 9276
rect 4704 9216 4768 9220
rect 4784 9276 4848 9280
rect 4784 9220 4788 9276
rect 4788 9220 4844 9276
rect 4844 9220 4848 9276
rect 4784 9216 4848 9220
rect 4864 9276 4928 9280
rect 4864 9220 4868 9276
rect 4868 9220 4924 9276
rect 4924 9220 4928 9276
rect 4864 9216 4928 9220
rect 7072 9276 7136 9280
rect 7072 9220 7076 9276
rect 7076 9220 7132 9276
rect 7132 9220 7136 9276
rect 7072 9216 7136 9220
rect 7152 9276 7216 9280
rect 7152 9220 7156 9276
rect 7156 9220 7212 9276
rect 7212 9220 7216 9276
rect 7152 9216 7216 9220
rect 7232 9276 7296 9280
rect 7232 9220 7236 9276
rect 7236 9220 7292 9276
rect 7292 9220 7296 9276
rect 7232 9216 7296 9220
rect 7312 9276 7376 9280
rect 7312 9220 7316 9276
rect 7316 9220 7372 9276
rect 7372 9220 7376 9276
rect 7312 9216 7376 9220
rect 9520 9276 9584 9280
rect 9520 9220 9524 9276
rect 9524 9220 9580 9276
rect 9580 9220 9584 9276
rect 9520 9216 9584 9220
rect 9600 9276 9664 9280
rect 9600 9220 9604 9276
rect 9604 9220 9660 9276
rect 9660 9220 9664 9276
rect 9600 9216 9664 9220
rect 9680 9276 9744 9280
rect 9680 9220 9684 9276
rect 9684 9220 9740 9276
rect 9740 9220 9744 9276
rect 9680 9216 9744 9220
rect 9760 9276 9824 9280
rect 9760 9220 9764 9276
rect 9764 9220 9820 9276
rect 9820 9220 9824 9276
rect 9760 9216 9824 9220
rect 3400 8732 3464 8736
rect 3400 8676 3404 8732
rect 3404 8676 3460 8732
rect 3460 8676 3464 8732
rect 3400 8672 3464 8676
rect 3480 8732 3544 8736
rect 3480 8676 3484 8732
rect 3484 8676 3540 8732
rect 3540 8676 3544 8732
rect 3480 8672 3544 8676
rect 3560 8732 3624 8736
rect 3560 8676 3564 8732
rect 3564 8676 3620 8732
rect 3620 8676 3624 8732
rect 3560 8672 3624 8676
rect 3640 8732 3704 8736
rect 3640 8676 3644 8732
rect 3644 8676 3700 8732
rect 3700 8676 3704 8732
rect 3640 8672 3704 8676
rect 5848 8732 5912 8736
rect 5848 8676 5852 8732
rect 5852 8676 5908 8732
rect 5908 8676 5912 8732
rect 5848 8672 5912 8676
rect 5928 8732 5992 8736
rect 5928 8676 5932 8732
rect 5932 8676 5988 8732
rect 5988 8676 5992 8732
rect 5928 8672 5992 8676
rect 6008 8732 6072 8736
rect 6008 8676 6012 8732
rect 6012 8676 6068 8732
rect 6068 8676 6072 8732
rect 6008 8672 6072 8676
rect 6088 8732 6152 8736
rect 6088 8676 6092 8732
rect 6092 8676 6148 8732
rect 6148 8676 6152 8732
rect 6088 8672 6152 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 8536 8732 8600 8736
rect 8536 8676 8540 8732
rect 8540 8676 8596 8732
rect 8596 8676 8600 8732
rect 8536 8672 8600 8676
rect 2176 8188 2240 8192
rect 2176 8132 2180 8188
rect 2180 8132 2236 8188
rect 2236 8132 2240 8188
rect 2176 8128 2240 8132
rect 2256 8188 2320 8192
rect 2256 8132 2260 8188
rect 2260 8132 2316 8188
rect 2316 8132 2320 8188
rect 2256 8128 2320 8132
rect 2336 8188 2400 8192
rect 2336 8132 2340 8188
rect 2340 8132 2396 8188
rect 2396 8132 2400 8188
rect 2336 8128 2400 8132
rect 2416 8188 2480 8192
rect 2416 8132 2420 8188
rect 2420 8132 2476 8188
rect 2476 8132 2480 8188
rect 2416 8128 2480 8132
rect 4624 8188 4688 8192
rect 4624 8132 4628 8188
rect 4628 8132 4684 8188
rect 4684 8132 4688 8188
rect 4624 8128 4688 8132
rect 4704 8188 4768 8192
rect 4704 8132 4708 8188
rect 4708 8132 4764 8188
rect 4764 8132 4768 8188
rect 4704 8128 4768 8132
rect 4784 8188 4848 8192
rect 4784 8132 4788 8188
rect 4788 8132 4844 8188
rect 4844 8132 4848 8188
rect 4784 8128 4848 8132
rect 4864 8188 4928 8192
rect 4864 8132 4868 8188
rect 4868 8132 4924 8188
rect 4924 8132 4928 8188
rect 4864 8128 4928 8132
rect 7072 8188 7136 8192
rect 7072 8132 7076 8188
rect 7076 8132 7132 8188
rect 7132 8132 7136 8188
rect 7072 8128 7136 8132
rect 7152 8188 7216 8192
rect 7152 8132 7156 8188
rect 7156 8132 7212 8188
rect 7212 8132 7216 8188
rect 7152 8128 7216 8132
rect 7232 8188 7296 8192
rect 7232 8132 7236 8188
rect 7236 8132 7292 8188
rect 7292 8132 7296 8188
rect 7232 8128 7296 8132
rect 7312 8188 7376 8192
rect 7312 8132 7316 8188
rect 7316 8132 7372 8188
rect 7372 8132 7376 8188
rect 7312 8128 7376 8132
rect 9520 8188 9584 8192
rect 9520 8132 9524 8188
rect 9524 8132 9580 8188
rect 9580 8132 9584 8188
rect 9520 8128 9584 8132
rect 9600 8188 9664 8192
rect 9600 8132 9604 8188
rect 9604 8132 9660 8188
rect 9660 8132 9664 8188
rect 9600 8128 9664 8132
rect 9680 8188 9744 8192
rect 9680 8132 9684 8188
rect 9684 8132 9740 8188
rect 9740 8132 9744 8188
rect 9680 8128 9744 8132
rect 9760 8188 9824 8192
rect 9760 8132 9764 8188
rect 9764 8132 9820 8188
rect 9820 8132 9824 8188
rect 9760 8128 9824 8132
rect 3400 7644 3464 7648
rect 3400 7588 3404 7644
rect 3404 7588 3460 7644
rect 3460 7588 3464 7644
rect 3400 7584 3464 7588
rect 3480 7644 3544 7648
rect 3480 7588 3484 7644
rect 3484 7588 3540 7644
rect 3540 7588 3544 7644
rect 3480 7584 3544 7588
rect 3560 7644 3624 7648
rect 3560 7588 3564 7644
rect 3564 7588 3620 7644
rect 3620 7588 3624 7644
rect 3560 7584 3624 7588
rect 3640 7644 3704 7648
rect 3640 7588 3644 7644
rect 3644 7588 3700 7644
rect 3700 7588 3704 7644
rect 3640 7584 3704 7588
rect 5848 7644 5912 7648
rect 5848 7588 5852 7644
rect 5852 7588 5908 7644
rect 5908 7588 5912 7644
rect 5848 7584 5912 7588
rect 5928 7644 5992 7648
rect 5928 7588 5932 7644
rect 5932 7588 5988 7644
rect 5988 7588 5992 7644
rect 5928 7584 5992 7588
rect 6008 7644 6072 7648
rect 6008 7588 6012 7644
rect 6012 7588 6068 7644
rect 6068 7588 6072 7644
rect 6008 7584 6072 7588
rect 6088 7644 6152 7648
rect 6088 7588 6092 7644
rect 6092 7588 6148 7644
rect 6148 7588 6152 7644
rect 6088 7584 6152 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 8536 7644 8600 7648
rect 8536 7588 8540 7644
rect 8540 7588 8596 7644
rect 8596 7588 8600 7644
rect 8536 7584 8600 7588
rect 2176 7100 2240 7104
rect 2176 7044 2180 7100
rect 2180 7044 2236 7100
rect 2236 7044 2240 7100
rect 2176 7040 2240 7044
rect 2256 7100 2320 7104
rect 2256 7044 2260 7100
rect 2260 7044 2316 7100
rect 2316 7044 2320 7100
rect 2256 7040 2320 7044
rect 2336 7100 2400 7104
rect 2336 7044 2340 7100
rect 2340 7044 2396 7100
rect 2396 7044 2400 7100
rect 2336 7040 2400 7044
rect 2416 7100 2480 7104
rect 2416 7044 2420 7100
rect 2420 7044 2476 7100
rect 2476 7044 2480 7100
rect 2416 7040 2480 7044
rect 4624 7100 4688 7104
rect 4624 7044 4628 7100
rect 4628 7044 4684 7100
rect 4684 7044 4688 7100
rect 4624 7040 4688 7044
rect 4704 7100 4768 7104
rect 4704 7044 4708 7100
rect 4708 7044 4764 7100
rect 4764 7044 4768 7100
rect 4704 7040 4768 7044
rect 4784 7100 4848 7104
rect 4784 7044 4788 7100
rect 4788 7044 4844 7100
rect 4844 7044 4848 7100
rect 4784 7040 4848 7044
rect 4864 7100 4928 7104
rect 4864 7044 4868 7100
rect 4868 7044 4924 7100
rect 4924 7044 4928 7100
rect 4864 7040 4928 7044
rect 7072 7100 7136 7104
rect 7072 7044 7076 7100
rect 7076 7044 7132 7100
rect 7132 7044 7136 7100
rect 7072 7040 7136 7044
rect 7152 7100 7216 7104
rect 7152 7044 7156 7100
rect 7156 7044 7212 7100
rect 7212 7044 7216 7100
rect 7152 7040 7216 7044
rect 7232 7100 7296 7104
rect 7232 7044 7236 7100
rect 7236 7044 7292 7100
rect 7292 7044 7296 7100
rect 7232 7040 7296 7044
rect 7312 7100 7376 7104
rect 7312 7044 7316 7100
rect 7316 7044 7372 7100
rect 7372 7044 7376 7100
rect 7312 7040 7376 7044
rect 9520 7100 9584 7104
rect 9520 7044 9524 7100
rect 9524 7044 9580 7100
rect 9580 7044 9584 7100
rect 9520 7040 9584 7044
rect 9600 7100 9664 7104
rect 9600 7044 9604 7100
rect 9604 7044 9660 7100
rect 9660 7044 9664 7100
rect 9600 7040 9664 7044
rect 9680 7100 9744 7104
rect 9680 7044 9684 7100
rect 9684 7044 9740 7100
rect 9740 7044 9744 7100
rect 9680 7040 9744 7044
rect 9760 7100 9824 7104
rect 9760 7044 9764 7100
rect 9764 7044 9820 7100
rect 9820 7044 9824 7100
rect 9760 7040 9824 7044
rect 3400 6556 3464 6560
rect 3400 6500 3404 6556
rect 3404 6500 3460 6556
rect 3460 6500 3464 6556
rect 3400 6496 3464 6500
rect 3480 6556 3544 6560
rect 3480 6500 3484 6556
rect 3484 6500 3540 6556
rect 3540 6500 3544 6556
rect 3480 6496 3544 6500
rect 3560 6556 3624 6560
rect 3560 6500 3564 6556
rect 3564 6500 3620 6556
rect 3620 6500 3624 6556
rect 3560 6496 3624 6500
rect 3640 6556 3704 6560
rect 3640 6500 3644 6556
rect 3644 6500 3700 6556
rect 3700 6500 3704 6556
rect 3640 6496 3704 6500
rect 5848 6556 5912 6560
rect 5848 6500 5852 6556
rect 5852 6500 5908 6556
rect 5908 6500 5912 6556
rect 5848 6496 5912 6500
rect 5928 6556 5992 6560
rect 5928 6500 5932 6556
rect 5932 6500 5988 6556
rect 5988 6500 5992 6556
rect 5928 6496 5992 6500
rect 6008 6556 6072 6560
rect 6008 6500 6012 6556
rect 6012 6500 6068 6556
rect 6068 6500 6072 6556
rect 6008 6496 6072 6500
rect 6088 6556 6152 6560
rect 6088 6500 6092 6556
rect 6092 6500 6148 6556
rect 6148 6500 6152 6556
rect 6088 6496 6152 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 8536 6556 8600 6560
rect 8536 6500 8540 6556
rect 8540 6500 8596 6556
rect 8596 6500 8600 6556
rect 8536 6496 8600 6500
rect 2176 6012 2240 6016
rect 2176 5956 2180 6012
rect 2180 5956 2236 6012
rect 2236 5956 2240 6012
rect 2176 5952 2240 5956
rect 2256 6012 2320 6016
rect 2256 5956 2260 6012
rect 2260 5956 2316 6012
rect 2316 5956 2320 6012
rect 2256 5952 2320 5956
rect 2336 6012 2400 6016
rect 2336 5956 2340 6012
rect 2340 5956 2396 6012
rect 2396 5956 2400 6012
rect 2336 5952 2400 5956
rect 2416 6012 2480 6016
rect 2416 5956 2420 6012
rect 2420 5956 2476 6012
rect 2476 5956 2480 6012
rect 2416 5952 2480 5956
rect 4624 6012 4688 6016
rect 4624 5956 4628 6012
rect 4628 5956 4684 6012
rect 4684 5956 4688 6012
rect 4624 5952 4688 5956
rect 4704 6012 4768 6016
rect 4704 5956 4708 6012
rect 4708 5956 4764 6012
rect 4764 5956 4768 6012
rect 4704 5952 4768 5956
rect 4784 6012 4848 6016
rect 4784 5956 4788 6012
rect 4788 5956 4844 6012
rect 4844 5956 4848 6012
rect 4784 5952 4848 5956
rect 4864 6012 4928 6016
rect 4864 5956 4868 6012
rect 4868 5956 4924 6012
rect 4924 5956 4928 6012
rect 4864 5952 4928 5956
rect 7072 6012 7136 6016
rect 7072 5956 7076 6012
rect 7076 5956 7132 6012
rect 7132 5956 7136 6012
rect 7072 5952 7136 5956
rect 7152 6012 7216 6016
rect 7152 5956 7156 6012
rect 7156 5956 7212 6012
rect 7212 5956 7216 6012
rect 7152 5952 7216 5956
rect 7232 6012 7296 6016
rect 7232 5956 7236 6012
rect 7236 5956 7292 6012
rect 7292 5956 7296 6012
rect 7232 5952 7296 5956
rect 7312 6012 7376 6016
rect 7312 5956 7316 6012
rect 7316 5956 7372 6012
rect 7372 5956 7376 6012
rect 7312 5952 7376 5956
rect 9520 6012 9584 6016
rect 9520 5956 9524 6012
rect 9524 5956 9580 6012
rect 9580 5956 9584 6012
rect 9520 5952 9584 5956
rect 9600 6012 9664 6016
rect 9600 5956 9604 6012
rect 9604 5956 9660 6012
rect 9660 5956 9664 6012
rect 9600 5952 9664 5956
rect 9680 6012 9744 6016
rect 9680 5956 9684 6012
rect 9684 5956 9740 6012
rect 9740 5956 9744 6012
rect 9680 5952 9744 5956
rect 9760 6012 9824 6016
rect 9760 5956 9764 6012
rect 9764 5956 9820 6012
rect 9820 5956 9824 6012
rect 9760 5952 9824 5956
rect 3400 5468 3464 5472
rect 3400 5412 3404 5468
rect 3404 5412 3460 5468
rect 3460 5412 3464 5468
rect 3400 5408 3464 5412
rect 3480 5468 3544 5472
rect 3480 5412 3484 5468
rect 3484 5412 3540 5468
rect 3540 5412 3544 5468
rect 3480 5408 3544 5412
rect 3560 5468 3624 5472
rect 3560 5412 3564 5468
rect 3564 5412 3620 5468
rect 3620 5412 3624 5468
rect 3560 5408 3624 5412
rect 3640 5468 3704 5472
rect 3640 5412 3644 5468
rect 3644 5412 3700 5468
rect 3700 5412 3704 5468
rect 3640 5408 3704 5412
rect 5848 5468 5912 5472
rect 5848 5412 5852 5468
rect 5852 5412 5908 5468
rect 5908 5412 5912 5468
rect 5848 5408 5912 5412
rect 5928 5468 5992 5472
rect 5928 5412 5932 5468
rect 5932 5412 5988 5468
rect 5988 5412 5992 5468
rect 5928 5408 5992 5412
rect 6008 5468 6072 5472
rect 6008 5412 6012 5468
rect 6012 5412 6068 5468
rect 6068 5412 6072 5468
rect 6008 5408 6072 5412
rect 6088 5468 6152 5472
rect 6088 5412 6092 5468
rect 6092 5412 6148 5468
rect 6148 5412 6152 5468
rect 6088 5408 6152 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 8536 5468 8600 5472
rect 8536 5412 8540 5468
rect 8540 5412 8596 5468
rect 8596 5412 8600 5468
rect 8536 5408 8600 5412
rect 2176 4924 2240 4928
rect 2176 4868 2180 4924
rect 2180 4868 2236 4924
rect 2236 4868 2240 4924
rect 2176 4864 2240 4868
rect 2256 4924 2320 4928
rect 2256 4868 2260 4924
rect 2260 4868 2316 4924
rect 2316 4868 2320 4924
rect 2256 4864 2320 4868
rect 2336 4924 2400 4928
rect 2336 4868 2340 4924
rect 2340 4868 2396 4924
rect 2396 4868 2400 4924
rect 2336 4864 2400 4868
rect 2416 4924 2480 4928
rect 2416 4868 2420 4924
rect 2420 4868 2476 4924
rect 2476 4868 2480 4924
rect 2416 4864 2480 4868
rect 4624 4924 4688 4928
rect 4624 4868 4628 4924
rect 4628 4868 4684 4924
rect 4684 4868 4688 4924
rect 4624 4864 4688 4868
rect 4704 4924 4768 4928
rect 4704 4868 4708 4924
rect 4708 4868 4764 4924
rect 4764 4868 4768 4924
rect 4704 4864 4768 4868
rect 4784 4924 4848 4928
rect 4784 4868 4788 4924
rect 4788 4868 4844 4924
rect 4844 4868 4848 4924
rect 4784 4864 4848 4868
rect 4864 4924 4928 4928
rect 4864 4868 4868 4924
rect 4868 4868 4924 4924
rect 4924 4868 4928 4924
rect 4864 4864 4928 4868
rect 7072 4924 7136 4928
rect 7072 4868 7076 4924
rect 7076 4868 7132 4924
rect 7132 4868 7136 4924
rect 7072 4864 7136 4868
rect 7152 4924 7216 4928
rect 7152 4868 7156 4924
rect 7156 4868 7212 4924
rect 7212 4868 7216 4924
rect 7152 4864 7216 4868
rect 7232 4924 7296 4928
rect 7232 4868 7236 4924
rect 7236 4868 7292 4924
rect 7292 4868 7296 4924
rect 7232 4864 7296 4868
rect 7312 4924 7376 4928
rect 7312 4868 7316 4924
rect 7316 4868 7372 4924
rect 7372 4868 7376 4924
rect 7312 4864 7376 4868
rect 9520 4924 9584 4928
rect 9520 4868 9524 4924
rect 9524 4868 9580 4924
rect 9580 4868 9584 4924
rect 9520 4864 9584 4868
rect 9600 4924 9664 4928
rect 9600 4868 9604 4924
rect 9604 4868 9660 4924
rect 9660 4868 9664 4924
rect 9600 4864 9664 4868
rect 9680 4924 9744 4928
rect 9680 4868 9684 4924
rect 9684 4868 9740 4924
rect 9740 4868 9744 4924
rect 9680 4864 9744 4868
rect 9760 4924 9824 4928
rect 9760 4868 9764 4924
rect 9764 4868 9820 4924
rect 9820 4868 9824 4924
rect 9760 4864 9824 4868
rect 3400 4380 3464 4384
rect 3400 4324 3404 4380
rect 3404 4324 3460 4380
rect 3460 4324 3464 4380
rect 3400 4320 3464 4324
rect 3480 4380 3544 4384
rect 3480 4324 3484 4380
rect 3484 4324 3540 4380
rect 3540 4324 3544 4380
rect 3480 4320 3544 4324
rect 3560 4380 3624 4384
rect 3560 4324 3564 4380
rect 3564 4324 3620 4380
rect 3620 4324 3624 4380
rect 3560 4320 3624 4324
rect 3640 4380 3704 4384
rect 3640 4324 3644 4380
rect 3644 4324 3700 4380
rect 3700 4324 3704 4380
rect 3640 4320 3704 4324
rect 5848 4380 5912 4384
rect 5848 4324 5852 4380
rect 5852 4324 5908 4380
rect 5908 4324 5912 4380
rect 5848 4320 5912 4324
rect 5928 4380 5992 4384
rect 5928 4324 5932 4380
rect 5932 4324 5988 4380
rect 5988 4324 5992 4380
rect 5928 4320 5992 4324
rect 6008 4380 6072 4384
rect 6008 4324 6012 4380
rect 6012 4324 6068 4380
rect 6068 4324 6072 4380
rect 6008 4320 6072 4324
rect 6088 4380 6152 4384
rect 6088 4324 6092 4380
rect 6092 4324 6148 4380
rect 6148 4324 6152 4380
rect 6088 4320 6152 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 8536 4380 8600 4384
rect 8536 4324 8540 4380
rect 8540 4324 8596 4380
rect 8596 4324 8600 4380
rect 8536 4320 8600 4324
rect 2176 3836 2240 3840
rect 2176 3780 2180 3836
rect 2180 3780 2236 3836
rect 2236 3780 2240 3836
rect 2176 3776 2240 3780
rect 2256 3836 2320 3840
rect 2256 3780 2260 3836
rect 2260 3780 2316 3836
rect 2316 3780 2320 3836
rect 2256 3776 2320 3780
rect 2336 3836 2400 3840
rect 2336 3780 2340 3836
rect 2340 3780 2396 3836
rect 2396 3780 2400 3836
rect 2336 3776 2400 3780
rect 2416 3836 2480 3840
rect 2416 3780 2420 3836
rect 2420 3780 2476 3836
rect 2476 3780 2480 3836
rect 2416 3776 2480 3780
rect 4624 3836 4688 3840
rect 4624 3780 4628 3836
rect 4628 3780 4684 3836
rect 4684 3780 4688 3836
rect 4624 3776 4688 3780
rect 4704 3836 4768 3840
rect 4704 3780 4708 3836
rect 4708 3780 4764 3836
rect 4764 3780 4768 3836
rect 4704 3776 4768 3780
rect 4784 3836 4848 3840
rect 4784 3780 4788 3836
rect 4788 3780 4844 3836
rect 4844 3780 4848 3836
rect 4784 3776 4848 3780
rect 4864 3836 4928 3840
rect 4864 3780 4868 3836
rect 4868 3780 4924 3836
rect 4924 3780 4928 3836
rect 4864 3776 4928 3780
rect 7072 3836 7136 3840
rect 7072 3780 7076 3836
rect 7076 3780 7132 3836
rect 7132 3780 7136 3836
rect 7072 3776 7136 3780
rect 7152 3836 7216 3840
rect 7152 3780 7156 3836
rect 7156 3780 7212 3836
rect 7212 3780 7216 3836
rect 7152 3776 7216 3780
rect 7232 3836 7296 3840
rect 7232 3780 7236 3836
rect 7236 3780 7292 3836
rect 7292 3780 7296 3836
rect 7232 3776 7296 3780
rect 7312 3836 7376 3840
rect 7312 3780 7316 3836
rect 7316 3780 7372 3836
rect 7372 3780 7376 3836
rect 7312 3776 7376 3780
rect 9520 3836 9584 3840
rect 9520 3780 9524 3836
rect 9524 3780 9580 3836
rect 9580 3780 9584 3836
rect 9520 3776 9584 3780
rect 9600 3836 9664 3840
rect 9600 3780 9604 3836
rect 9604 3780 9660 3836
rect 9660 3780 9664 3836
rect 9600 3776 9664 3780
rect 9680 3836 9744 3840
rect 9680 3780 9684 3836
rect 9684 3780 9740 3836
rect 9740 3780 9744 3836
rect 9680 3776 9744 3780
rect 9760 3836 9824 3840
rect 9760 3780 9764 3836
rect 9764 3780 9820 3836
rect 9820 3780 9824 3836
rect 9760 3776 9824 3780
rect 3400 3292 3464 3296
rect 3400 3236 3404 3292
rect 3404 3236 3460 3292
rect 3460 3236 3464 3292
rect 3400 3232 3464 3236
rect 3480 3292 3544 3296
rect 3480 3236 3484 3292
rect 3484 3236 3540 3292
rect 3540 3236 3544 3292
rect 3480 3232 3544 3236
rect 3560 3292 3624 3296
rect 3560 3236 3564 3292
rect 3564 3236 3620 3292
rect 3620 3236 3624 3292
rect 3560 3232 3624 3236
rect 3640 3292 3704 3296
rect 3640 3236 3644 3292
rect 3644 3236 3700 3292
rect 3700 3236 3704 3292
rect 3640 3232 3704 3236
rect 5848 3292 5912 3296
rect 5848 3236 5852 3292
rect 5852 3236 5908 3292
rect 5908 3236 5912 3292
rect 5848 3232 5912 3236
rect 5928 3292 5992 3296
rect 5928 3236 5932 3292
rect 5932 3236 5988 3292
rect 5988 3236 5992 3292
rect 5928 3232 5992 3236
rect 6008 3292 6072 3296
rect 6008 3236 6012 3292
rect 6012 3236 6068 3292
rect 6068 3236 6072 3292
rect 6008 3232 6072 3236
rect 6088 3292 6152 3296
rect 6088 3236 6092 3292
rect 6092 3236 6148 3292
rect 6148 3236 6152 3292
rect 6088 3232 6152 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 8536 3292 8600 3296
rect 8536 3236 8540 3292
rect 8540 3236 8596 3292
rect 8596 3236 8600 3292
rect 8536 3232 8600 3236
rect 2176 2748 2240 2752
rect 2176 2692 2180 2748
rect 2180 2692 2236 2748
rect 2236 2692 2240 2748
rect 2176 2688 2240 2692
rect 2256 2748 2320 2752
rect 2256 2692 2260 2748
rect 2260 2692 2316 2748
rect 2316 2692 2320 2748
rect 2256 2688 2320 2692
rect 2336 2748 2400 2752
rect 2336 2692 2340 2748
rect 2340 2692 2396 2748
rect 2396 2692 2400 2748
rect 2336 2688 2400 2692
rect 2416 2748 2480 2752
rect 2416 2692 2420 2748
rect 2420 2692 2476 2748
rect 2476 2692 2480 2748
rect 2416 2688 2480 2692
rect 4624 2748 4688 2752
rect 4624 2692 4628 2748
rect 4628 2692 4684 2748
rect 4684 2692 4688 2748
rect 4624 2688 4688 2692
rect 4704 2748 4768 2752
rect 4704 2692 4708 2748
rect 4708 2692 4764 2748
rect 4764 2692 4768 2748
rect 4704 2688 4768 2692
rect 4784 2748 4848 2752
rect 4784 2692 4788 2748
rect 4788 2692 4844 2748
rect 4844 2692 4848 2748
rect 4784 2688 4848 2692
rect 4864 2748 4928 2752
rect 4864 2692 4868 2748
rect 4868 2692 4924 2748
rect 4924 2692 4928 2748
rect 4864 2688 4928 2692
rect 7072 2748 7136 2752
rect 7072 2692 7076 2748
rect 7076 2692 7132 2748
rect 7132 2692 7136 2748
rect 7072 2688 7136 2692
rect 7152 2748 7216 2752
rect 7152 2692 7156 2748
rect 7156 2692 7212 2748
rect 7212 2692 7216 2748
rect 7152 2688 7216 2692
rect 7232 2748 7296 2752
rect 7232 2692 7236 2748
rect 7236 2692 7292 2748
rect 7292 2692 7296 2748
rect 7232 2688 7296 2692
rect 7312 2748 7376 2752
rect 7312 2692 7316 2748
rect 7316 2692 7372 2748
rect 7372 2692 7376 2748
rect 7312 2688 7376 2692
rect 9520 2748 9584 2752
rect 9520 2692 9524 2748
rect 9524 2692 9580 2748
rect 9580 2692 9584 2748
rect 9520 2688 9584 2692
rect 9600 2748 9664 2752
rect 9600 2692 9604 2748
rect 9604 2692 9660 2748
rect 9660 2692 9664 2748
rect 9600 2688 9664 2692
rect 9680 2748 9744 2752
rect 9680 2692 9684 2748
rect 9684 2692 9740 2748
rect 9740 2692 9744 2748
rect 9680 2688 9744 2692
rect 9760 2748 9824 2752
rect 9760 2692 9764 2748
rect 9764 2692 9820 2748
rect 9820 2692 9824 2748
rect 9760 2688 9824 2692
rect 3400 2204 3464 2208
rect 3400 2148 3404 2204
rect 3404 2148 3460 2204
rect 3460 2148 3464 2204
rect 3400 2144 3464 2148
rect 3480 2204 3544 2208
rect 3480 2148 3484 2204
rect 3484 2148 3540 2204
rect 3540 2148 3544 2204
rect 3480 2144 3544 2148
rect 3560 2204 3624 2208
rect 3560 2148 3564 2204
rect 3564 2148 3620 2204
rect 3620 2148 3624 2204
rect 3560 2144 3624 2148
rect 3640 2204 3704 2208
rect 3640 2148 3644 2204
rect 3644 2148 3700 2204
rect 3700 2148 3704 2204
rect 3640 2144 3704 2148
rect 5848 2204 5912 2208
rect 5848 2148 5852 2204
rect 5852 2148 5908 2204
rect 5908 2148 5912 2204
rect 5848 2144 5912 2148
rect 5928 2204 5992 2208
rect 5928 2148 5932 2204
rect 5932 2148 5988 2204
rect 5988 2148 5992 2204
rect 5928 2144 5992 2148
rect 6008 2204 6072 2208
rect 6008 2148 6012 2204
rect 6012 2148 6068 2204
rect 6068 2148 6072 2204
rect 6008 2144 6072 2148
rect 6088 2204 6152 2208
rect 6088 2148 6092 2204
rect 6092 2148 6148 2204
rect 6148 2148 6152 2204
rect 6088 2144 6152 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 8536 2204 8600 2208
rect 8536 2148 8540 2204
rect 8540 2148 8596 2204
rect 8596 2148 8600 2204
rect 8536 2144 8600 2148
<< metal4 >>
rect 2168 11456 2488 11472
rect 2168 11392 2176 11456
rect 2240 11392 2256 11456
rect 2320 11392 2336 11456
rect 2400 11392 2416 11456
rect 2480 11392 2488 11456
rect 2168 10368 2488 11392
rect 2168 10304 2176 10368
rect 2240 10304 2256 10368
rect 2320 10304 2336 10368
rect 2400 10304 2416 10368
rect 2480 10304 2488 10368
rect 2168 9280 2488 10304
rect 2168 9216 2176 9280
rect 2240 9216 2256 9280
rect 2320 9216 2336 9280
rect 2400 9216 2416 9280
rect 2480 9216 2488 9280
rect 2168 8192 2488 9216
rect 2168 8128 2176 8192
rect 2240 8128 2256 8192
rect 2320 8128 2336 8192
rect 2400 8128 2416 8192
rect 2480 8128 2488 8192
rect 2168 7104 2488 8128
rect 2168 7040 2176 7104
rect 2240 7040 2256 7104
rect 2320 7040 2336 7104
rect 2400 7040 2416 7104
rect 2480 7040 2488 7104
rect 2168 6016 2488 7040
rect 2168 5952 2176 6016
rect 2240 5952 2256 6016
rect 2320 5952 2336 6016
rect 2400 5952 2416 6016
rect 2480 5952 2488 6016
rect 2168 4928 2488 5952
rect 2168 4864 2176 4928
rect 2240 4864 2256 4928
rect 2320 4864 2336 4928
rect 2400 4864 2416 4928
rect 2480 4864 2488 4928
rect 2168 3840 2488 4864
rect 2168 3776 2176 3840
rect 2240 3776 2256 3840
rect 2320 3776 2336 3840
rect 2400 3776 2416 3840
rect 2480 3776 2488 3840
rect 2168 2752 2488 3776
rect 2168 2688 2176 2752
rect 2240 2688 2256 2752
rect 2320 2688 2336 2752
rect 2400 2688 2416 2752
rect 2480 2688 2488 2752
rect 2168 2128 2488 2688
rect 3392 10912 3712 11472
rect 3392 10848 3400 10912
rect 3464 10848 3480 10912
rect 3544 10848 3560 10912
rect 3624 10848 3640 10912
rect 3704 10848 3712 10912
rect 3392 9824 3712 10848
rect 3392 9760 3400 9824
rect 3464 9760 3480 9824
rect 3544 9760 3560 9824
rect 3624 9760 3640 9824
rect 3704 9760 3712 9824
rect 3392 8736 3712 9760
rect 3392 8672 3400 8736
rect 3464 8672 3480 8736
rect 3544 8672 3560 8736
rect 3624 8672 3640 8736
rect 3704 8672 3712 8736
rect 3392 7648 3712 8672
rect 3392 7584 3400 7648
rect 3464 7584 3480 7648
rect 3544 7584 3560 7648
rect 3624 7584 3640 7648
rect 3704 7584 3712 7648
rect 3392 6560 3712 7584
rect 3392 6496 3400 6560
rect 3464 6496 3480 6560
rect 3544 6496 3560 6560
rect 3624 6496 3640 6560
rect 3704 6496 3712 6560
rect 3392 5472 3712 6496
rect 3392 5408 3400 5472
rect 3464 5408 3480 5472
rect 3544 5408 3560 5472
rect 3624 5408 3640 5472
rect 3704 5408 3712 5472
rect 3392 4384 3712 5408
rect 3392 4320 3400 4384
rect 3464 4320 3480 4384
rect 3544 4320 3560 4384
rect 3624 4320 3640 4384
rect 3704 4320 3712 4384
rect 3392 3296 3712 4320
rect 3392 3232 3400 3296
rect 3464 3232 3480 3296
rect 3544 3232 3560 3296
rect 3624 3232 3640 3296
rect 3704 3232 3712 3296
rect 3392 2208 3712 3232
rect 3392 2144 3400 2208
rect 3464 2144 3480 2208
rect 3544 2144 3560 2208
rect 3624 2144 3640 2208
rect 3704 2144 3712 2208
rect 3392 2128 3712 2144
rect 4616 11456 4936 11472
rect 4616 11392 4624 11456
rect 4688 11392 4704 11456
rect 4768 11392 4784 11456
rect 4848 11392 4864 11456
rect 4928 11392 4936 11456
rect 4616 10368 4936 11392
rect 4616 10304 4624 10368
rect 4688 10304 4704 10368
rect 4768 10304 4784 10368
rect 4848 10304 4864 10368
rect 4928 10304 4936 10368
rect 4616 9280 4936 10304
rect 4616 9216 4624 9280
rect 4688 9216 4704 9280
rect 4768 9216 4784 9280
rect 4848 9216 4864 9280
rect 4928 9216 4936 9280
rect 4616 8192 4936 9216
rect 4616 8128 4624 8192
rect 4688 8128 4704 8192
rect 4768 8128 4784 8192
rect 4848 8128 4864 8192
rect 4928 8128 4936 8192
rect 4616 7104 4936 8128
rect 4616 7040 4624 7104
rect 4688 7040 4704 7104
rect 4768 7040 4784 7104
rect 4848 7040 4864 7104
rect 4928 7040 4936 7104
rect 4616 6016 4936 7040
rect 4616 5952 4624 6016
rect 4688 5952 4704 6016
rect 4768 5952 4784 6016
rect 4848 5952 4864 6016
rect 4928 5952 4936 6016
rect 4616 4928 4936 5952
rect 4616 4864 4624 4928
rect 4688 4864 4704 4928
rect 4768 4864 4784 4928
rect 4848 4864 4864 4928
rect 4928 4864 4936 4928
rect 4616 3840 4936 4864
rect 4616 3776 4624 3840
rect 4688 3776 4704 3840
rect 4768 3776 4784 3840
rect 4848 3776 4864 3840
rect 4928 3776 4936 3840
rect 4616 2752 4936 3776
rect 4616 2688 4624 2752
rect 4688 2688 4704 2752
rect 4768 2688 4784 2752
rect 4848 2688 4864 2752
rect 4928 2688 4936 2752
rect 4616 2128 4936 2688
rect 5840 10912 6160 11472
rect 5840 10848 5848 10912
rect 5912 10848 5928 10912
rect 5992 10848 6008 10912
rect 6072 10848 6088 10912
rect 6152 10848 6160 10912
rect 5840 9824 6160 10848
rect 5840 9760 5848 9824
rect 5912 9760 5928 9824
rect 5992 9760 6008 9824
rect 6072 9760 6088 9824
rect 6152 9760 6160 9824
rect 5840 8736 6160 9760
rect 5840 8672 5848 8736
rect 5912 8672 5928 8736
rect 5992 8672 6008 8736
rect 6072 8672 6088 8736
rect 6152 8672 6160 8736
rect 5840 7648 6160 8672
rect 5840 7584 5848 7648
rect 5912 7584 5928 7648
rect 5992 7584 6008 7648
rect 6072 7584 6088 7648
rect 6152 7584 6160 7648
rect 5840 6560 6160 7584
rect 5840 6496 5848 6560
rect 5912 6496 5928 6560
rect 5992 6496 6008 6560
rect 6072 6496 6088 6560
rect 6152 6496 6160 6560
rect 5840 5472 6160 6496
rect 5840 5408 5848 5472
rect 5912 5408 5928 5472
rect 5992 5408 6008 5472
rect 6072 5408 6088 5472
rect 6152 5408 6160 5472
rect 5840 4384 6160 5408
rect 5840 4320 5848 4384
rect 5912 4320 5928 4384
rect 5992 4320 6008 4384
rect 6072 4320 6088 4384
rect 6152 4320 6160 4384
rect 5840 3296 6160 4320
rect 5840 3232 5848 3296
rect 5912 3232 5928 3296
rect 5992 3232 6008 3296
rect 6072 3232 6088 3296
rect 6152 3232 6160 3296
rect 5840 2208 6160 3232
rect 5840 2144 5848 2208
rect 5912 2144 5928 2208
rect 5992 2144 6008 2208
rect 6072 2144 6088 2208
rect 6152 2144 6160 2208
rect 5840 2128 6160 2144
rect 7064 11456 7384 11472
rect 7064 11392 7072 11456
rect 7136 11392 7152 11456
rect 7216 11392 7232 11456
rect 7296 11392 7312 11456
rect 7376 11392 7384 11456
rect 7064 10368 7384 11392
rect 7064 10304 7072 10368
rect 7136 10304 7152 10368
rect 7216 10304 7232 10368
rect 7296 10304 7312 10368
rect 7376 10304 7384 10368
rect 7064 9280 7384 10304
rect 7064 9216 7072 9280
rect 7136 9216 7152 9280
rect 7216 9216 7232 9280
rect 7296 9216 7312 9280
rect 7376 9216 7384 9280
rect 7064 8192 7384 9216
rect 7064 8128 7072 8192
rect 7136 8128 7152 8192
rect 7216 8128 7232 8192
rect 7296 8128 7312 8192
rect 7376 8128 7384 8192
rect 7064 7104 7384 8128
rect 7064 7040 7072 7104
rect 7136 7040 7152 7104
rect 7216 7040 7232 7104
rect 7296 7040 7312 7104
rect 7376 7040 7384 7104
rect 7064 6016 7384 7040
rect 7064 5952 7072 6016
rect 7136 5952 7152 6016
rect 7216 5952 7232 6016
rect 7296 5952 7312 6016
rect 7376 5952 7384 6016
rect 7064 4928 7384 5952
rect 7064 4864 7072 4928
rect 7136 4864 7152 4928
rect 7216 4864 7232 4928
rect 7296 4864 7312 4928
rect 7376 4864 7384 4928
rect 7064 3840 7384 4864
rect 7064 3776 7072 3840
rect 7136 3776 7152 3840
rect 7216 3776 7232 3840
rect 7296 3776 7312 3840
rect 7376 3776 7384 3840
rect 7064 2752 7384 3776
rect 7064 2688 7072 2752
rect 7136 2688 7152 2752
rect 7216 2688 7232 2752
rect 7296 2688 7312 2752
rect 7376 2688 7384 2752
rect 7064 2128 7384 2688
rect 8288 10912 8608 11472
rect 8288 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8536 10912
rect 8600 10848 8608 10912
rect 8288 9824 8608 10848
rect 8288 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8536 9824
rect 8600 9760 8608 9824
rect 8288 8736 8608 9760
rect 8288 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8536 8736
rect 8600 8672 8608 8736
rect 8288 7648 8608 8672
rect 8288 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8536 7648
rect 8600 7584 8608 7648
rect 8288 6560 8608 7584
rect 8288 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8536 6560
rect 8600 6496 8608 6560
rect 8288 5472 8608 6496
rect 8288 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8536 5472
rect 8600 5408 8608 5472
rect 8288 4384 8608 5408
rect 8288 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8536 4384
rect 8600 4320 8608 4384
rect 8288 3296 8608 4320
rect 8288 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8536 3296
rect 8600 3232 8608 3296
rect 8288 2208 8608 3232
rect 8288 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8536 2208
rect 8600 2144 8608 2208
rect 8288 2128 8608 2144
rect 9512 11456 9832 11472
rect 9512 11392 9520 11456
rect 9584 11392 9600 11456
rect 9664 11392 9680 11456
rect 9744 11392 9760 11456
rect 9824 11392 9832 11456
rect 9512 10368 9832 11392
rect 9512 10304 9520 10368
rect 9584 10304 9600 10368
rect 9664 10304 9680 10368
rect 9744 10304 9760 10368
rect 9824 10304 9832 10368
rect 9512 9280 9832 10304
rect 9512 9216 9520 9280
rect 9584 9216 9600 9280
rect 9664 9216 9680 9280
rect 9744 9216 9760 9280
rect 9824 9216 9832 9280
rect 9512 8192 9832 9216
rect 9512 8128 9520 8192
rect 9584 8128 9600 8192
rect 9664 8128 9680 8192
rect 9744 8128 9760 8192
rect 9824 8128 9832 8192
rect 9512 7104 9832 8128
rect 9512 7040 9520 7104
rect 9584 7040 9600 7104
rect 9664 7040 9680 7104
rect 9744 7040 9760 7104
rect 9824 7040 9832 7104
rect 9512 6016 9832 7040
rect 9512 5952 9520 6016
rect 9584 5952 9600 6016
rect 9664 5952 9680 6016
rect 9744 5952 9760 6016
rect 9824 5952 9832 6016
rect 9512 4928 9832 5952
rect 9512 4864 9520 4928
rect 9584 4864 9600 4928
rect 9664 4864 9680 4928
rect 9744 4864 9760 4928
rect 9824 4864 9832 4928
rect 9512 3840 9832 4864
rect 9512 3776 9520 3840
rect 9584 3776 9600 3840
rect 9664 3776 9680 3840
rect 9744 3776 9760 3840
rect 9824 3776 9832 3840
rect 9512 2752 9832 3776
rect 9512 2688 9520 2752
rect 9584 2688 9600 2752
rect 9664 2688 9680 2752
rect 9744 2688 9760 2752
rect 9824 2688 9832 2752
rect 9512 2128 9832 2688
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_89
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1649977179
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_20
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_57
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  conb_1\[0\] dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[1\]
timestamp 1649977179
transform -1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[2\]
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[3\]
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[4\]
timestamp 1649977179
transform -1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[5\]
timestamp 1649977179
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[6\]
timestamp 1649977179
transform 1 0 9016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[7\]
timestamp 1649977179
transform 1 0 9016 0 1 4352
box -38 -48 314 592
<< labels >>
flabel metal4 s 3392 2128 3712 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5840 2128 6160 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8288 2128 8608 11472 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2168 2128 2488 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4616 2128 4936 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7064 2128 7384 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9512 2128 9832 11472 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 x[0]
port 2 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 x[1]
port 3 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 x[2]
port 4 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 x[3]
port 5 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 x[4]
port 6 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 x[5]
port 7 nsew signal tristate
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 x[6]
port 8 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 x[7]
port 9 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 12000 14000
<< end >>
