//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module const0
(
    const0
);

    output const0;

    wire \<const0> = 0 ;
    wire const0;

assign const0 = \<const0> ;
endmodule

