VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_tile
  CLASS BLOCK ;
  FOREIGN top_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 255.000 BY 285.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.720 10.640 91.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.720 10.640 141.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 10.640 191.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.720 10.640 241.320 272.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.720 10.640 16.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 10.640 116.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.720 10.640 166.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.720 10.640 216.320 272.240 ;
    END
  END VPWR
  PIN bottom_width_0_height_0_subtile_0__pin_cout_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_cout_0_
  PIN bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 16.190 281.000 16.470 285.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN bottom_width_0_height_0_subtile_0__pin_reg_out_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END bottom_width_0_height_0_subtile_0__pin_reg_out_0_
  PIN bottom_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 25.850 281.000 26.130 285.000 ;
    END
  END bottom_width_0_height_0_subtile_1__pin_inpad_0_
  PIN bottom_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 35.510 281.000 35.790 285.000 ;
    END
  END bottom_width_0_height_0_subtile_2__pin_inpad_0_
  PIN bottom_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 45.170 281.000 45.450 285.000 ;
    END
  END bottom_width_0_height_0_subtile_3__pin_inpad_0_
  PIN ccff_head_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END ccff_head_1
  PIN ccff_head_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 248.030 281.000 248.310 285.000 ;
    END
  END ccff_head_2
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 3.440 255.000 4.040 ;
    END
  END ccff_tail
  PIN ccff_tail_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 6.530 281.000 6.810 285.000 ;
    END
  END ccff_tail_0
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END chanx_left_in[29]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END chanx_left_out[29]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 129.920 255.000 130.520 ;
    END
  END chanx_right_in_0[0]
  PIN chanx_right_in_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 170.720 255.000 171.320 ;
    END
  END chanx_right_in_0[10]
  PIN chanx_right_in_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 174.800 255.000 175.400 ;
    END
  END chanx_right_in_0[11]
  PIN chanx_right_in_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 178.880 255.000 179.480 ;
    END
  END chanx_right_in_0[12]
  PIN chanx_right_in_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 182.960 255.000 183.560 ;
    END
  END chanx_right_in_0[13]
  PIN chanx_right_in_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 187.040 255.000 187.640 ;
    END
  END chanx_right_in_0[14]
  PIN chanx_right_in_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 191.120 255.000 191.720 ;
    END
  END chanx_right_in_0[15]
  PIN chanx_right_in_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 195.200 255.000 195.800 ;
    END
  END chanx_right_in_0[16]
  PIN chanx_right_in_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 199.280 255.000 199.880 ;
    END
  END chanx_right_in_0[17]
  PIN chanx_right_in_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 203.360 255.000 203.960 ;
    END
  END chanx_right_in_0[18]
  PIN chanx_right_in_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 207.440 255.000 208.040 ;
    END
  END chanx_right_in_0[19]
  PIN chanx_right_in_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 134.000 255.000 134.600 ;
    END
  END chanx_right_in_0[1]
  PIN chanx_right_in_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 211.520 255.000 212.120 ;
    END
  END chanx_right_in_0[20]
  PIN chanx_right_in_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 215.600 255.000 216.200 ;
    END
  END chanx_right_in_0[21]
  PIN chanx_right_in_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 219.680 255.000 220.280 ;
    END
  END chanx_right_in_0[22]
  PIN chanx_right_in_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 223.760 255.000 224.360 ;
    END
  END chanx_right_in_0[23]
  PIN chanx_right_in_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 227.840 255.000 228.440 ;
    END
  END chanx_right_in_0[24]
  PIN chanx_right_in_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 231.920 255.000 232.520 ;
    END
  END chanx_right_in_0[25]
  PIN chanx_right_in_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 236.000 255.000 236.600 ;
    END
  END chanx_right_in_0[26]
  PIN chanx_right_in_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 240.080 255.000 240.680 ;
    END
  END chanx_right_in_0[27]
  PIN chanx_right_in_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 244.160 255.000 244.760 ;
    END
  END chanx_right_in_0[28]
  PIN chanx_right_in_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 248.240 255.000 248.840 ;
    END
  END chanx_right_in_0[29]
  PIN chanx_right_in_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 138.080 255.000 138.680 ;
    END
  END chanx_right_in_0[2]
  PIN chanx_right_in_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 142.160 255.000 142.760 ;
    END
  END chanx_right_in_0[3]
  PIN chanx_right_in_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 146.240 255.000 146.840 ;
    END
  END chanx_right_in_0[4]
  PIN chanx_right_in_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 150.320 255.000 150.920 ;
    END
  END chanx_right_in_0[5]
  PIN chanx_right_in_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 154.400 255.000 155.000 ;
    END
  END chanx_right_in_0[6]
  PIN chanx_right_in_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 158.480 255.000 159.080 ;
    END
  END chanx_right_in_0[7]
  PIN chanx_right_in_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 162.560 255.000 163.160 ;
    END
  END chanx_right_in_0[8]
  PIN chanx_right_in_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 166.640 255.000 167.240 ;
    END
  END chanx_right_in_0[9]
  PIN chanx_right_out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 7.520 255.000 8.120 ;
    END
  END chanx_right_out_0[0]
  PIN chanx_right_out_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 48.320 255.000 48.920 ;
    END
  END chanx_right_out_0[10]
  PIN chanx_right_out_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 52.400 255.000 53.000 ;
    END
  END chanx_right_out_0[11]
  PIN chanx_right_out_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 56.480 255.000 57.080 ;
    END
  END chanx_right_out_0[12]
  PIN chanx_right_out_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 60.560 255.000 61.160 ;
    END
  END chanx_right_out_0[13]
  PIN chanx_right_out_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 64.640 255.000 65.240 ;
    END
  END chanx_right_out_0[14]
  PIN chanx_right_out_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 68.720 255.000 69.320 ;
    END
  END chanx_right_out_0[15]
  PIN chanx_right_out_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 72.800 255.000 73.400 ;
    END
  END chanx_right_out_0[16]
  PIN chanx_right_out_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 76.880 255.000 77.480 ;
    END
  END chanx_right_out_0[17]
  PIN chanx_right_out_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 80.960 255.000 81.560 ;
    END
  END chanx_right_out_0[18]
  PIN chanx_right_out_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 85.040 255.000 85.640 ;
    END
  END chanx_right_out_0[19]
  PIN chanx_right_out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 11.600 255.000 12.200 ;
    END
  END chanx_right_out_0[1]
  PIN chanx_right_out_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 89.120 255.000 89.720 ;
    END
  END chanx_right_out_0[20]
  PIN chanx_right_out_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 93.200 255.000 93.800 ;
    END
  END chanx_right_out_0[21]
  PIN chanx_right_out_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 97.280 255.000 97.880 ;
    END
  END chanx_right_out_0[22]
  PIN chanx_right_out_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 101.360 255.000 101.960 ;
    END
  END chanx_right_out_0[23]
  PIN chanx_right_out_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 105.440 255.000 106.040 ;
    END
  END chanx_right_out_0[24]
  PIN chanx_right_out_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 109.520 255.000 110.120 ;
    END
  END chanx_right_out_0[25]
  PIN chanx_right_out_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 113.600 255.000 114.200 ;
    END
  END chanx_right_out_0[26]
  PIN chanx_right_out_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 117.680 255.000 118.280 ;
    END
  END chanx_right_out_0[27]
  PIN chanx_right_out_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 121.760 255.000 122.360 ;
    END
  END chanx_right_out_0[28]
  PIN chanx_right_out_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 125.840 255.000 126.440 ;
    END
  END chanx_right_out_0[29]
  PIN chanx_right_out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 15.680 255.000 16.280 ;
    END
  END chanx_right_out_0[2]
  PIN chanx_right_out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 19.760 255.000 20.360 ;
    END
  END chanx_right_out_0[3]
  PIN chanx_right_out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 23.840 255.000 24.440 ;
    END
  END chanx_right_out_0[4]
  PIN chanx_right_out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 27.920 255.000 28.520 ;
    END
  END chanx_right_out_0[5]
  PIN chanx_right_out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 32.000 255.000 32.600 ;
    END
  END chanx_right_out_0[6]
  PIN chanx_right_out_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 36.080 255.000 36.680 ;
    END
  END chanx_right_out_0[7]
  PIN chanx_right_out_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 40.160 255.000 40.760 ;
    END
  END chanx_right_out_0[8]
  PIN chanx_right_out_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 251.000 44.240 255.000 44.840 ;
    END
  END chanx_right_out_0[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END chany_bottom_in[29]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END chany_bottom_out[29]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END chany_bottom_out[9]
  PIN clk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END clk0
  PIN gfpga_pad_io_soc_dir[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 54.830 281.000 55.110 285.000 ;
    END
  END gfpga_pad_io_soc_dir[0]
  PIN gfpga_pad_io_soc_dir[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 64.490 281.000 64.770 285.000 ;
    END
  END gfpga_pad_io_soc_dir[1]
  PIN gfpga_pad_io_soc_dir[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 74.150 281.000 74.430 285.000 ;
    END
  END gfpga_pad_io_soc_dir[2]
  PIN gfpga_pad_io_soc_dir[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 83.810 281.000 84.090 285.000 ;
    END
  END gfpga_pad_io_soc_dir[3]
  PIN gfpga_pad_io_soc_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 281.000 132.390 285.000 ;
    END
  END gfpga_pad_io_soc_in[0]
  PIN gfpga_pad_io_soc_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 281.000 142.050 285.000 ;
    END
  END gfpga_pad_io_soc_in[1]
  PIN gfpga_pad_io_soc_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 281.000 151.710 285.000 ;
    END
  END gfpga_pad_io_soc_in[2]
  PIN gfpga_pad_io_soc_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 281.000 161.370 285.000 ;
    END
  END gfpga_pad_io_soc_in[3]
  PIN gfpga_pad_io_soc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 93.470 281.000 93.750 285.000 ;
    END
  END gfpga_pad_io_soc_out[0]
  PIN gfpga_pad_io_soc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 103.130 281.000 103.410 285.000 ;
    END
  END gfpga_pad_io_soc_out[1]
  PIN gfpga_pad_io_soc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 112.790 281.000 113.070 285.000 ;
    END
  END gfpga_pad_io_soc_out[2]
  PIN gfpga_pad_io_soc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 122.450 281.000 122.730 285.000 ;
    END
  END gfpga_pad_io_soc_out[3]
  PIN isol_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 281.000 171.030 285.000 ;
    END
  END isol_n
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END prog_clk
  PIN prog_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END prog_reset
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END reset
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 252.320 255.000 252.920 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 256.400 255.000 257.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 260.480 255.000 261.080 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 264.560 255.000 265.160 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 268.640 255.000 269.240 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 272.720 255.000 273.320 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 276.800 255.000 277.400 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met3 ;
        RECT 251.000 280.880 255.000 281.480 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 281.000 180.690 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 190.070 281.000 190.350 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 281.000 200.010 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 281.000 209.670 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
  PIN right_width_0_height_0_subtile_0__pin_O_10_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_10_
  PIN right_width_0_height_0_subtile_0__pin_O_11_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_11_
  PIN right_width_0_height_0_subtile_0__pin_O_12_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_12_
  PIN right_width_0_height_0_subtile_0__pin_O_13_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_13_
  PIN right_width_0_height_0_subtile_0__pin_O_14_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_14_
  PIN right_width_0_height_0_subtile_0__pin_O_15_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_15_
  PIN right_width_0_height_0_subtile_0__pin_O_8_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_8_
  PIN right_width_0_height_0_subtile_0__pin_O_9_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END right_width_0_height_0_subtile_0__pin_O_9_
  PIN sc_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 281.000 238.650 285.000 ;
    END
  END sc_in
  PIN sc_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END sc_out
  PIN test_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END test_enable
  PIN top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_0_
  PIN top_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_1_
  PIN top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_2_
  PIN top_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_3_
  PIN top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_4_
  PIN top_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_5_
  PIN top_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_6_
  PIN top_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END top_width_0_height_0_subtile_0__pin_O_7_
  PIN top_width_0_height_0_subtile_0__pin_cin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 281.000 219.330 285.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_cin_0_
  PIN top_width_0_height_0_subtile_0__pin_reg_in_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.110000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 281.000 228.990 285.000 ;
    END
  END top_width_0_height_0_subtile_0__pin_reg_in_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 249.320 272.085 ;
      LAYER met1 ;
        RECT 3.290 8.200 249.320 272.640 ;
      LAYER met2 ;
        RECT 3.320 280.720 6.250 281.365 ;
        RECT 7.090 280.720 15.910 281.365 ;
        RECT 16.750 280.720 25.570 281.365 ;
        RECT 26.410 280.720 35.230 281.365 ;
        RECT 36.070 280.720 44.890 281.365 ;
        RECT 45.730 280.720 54.550 281.365 ;
        RECT 55.390 280.720 64.210 281.365 ;
        RECT 65.050 280.720 73.870 281.365 ;
        RECT 74.710 280.720 83.530 281.365 ;
        RECT 84.370 280.720 93.190 281.365 ;
        RECT 94.030 280.720 102.850 281.365 ;
        RECT 103.690 280.720 112.510 281.365 ;
        RECT 113.350 280.720 122.170 281.365 ;
        RECT 123.010 280.720 131.830 281.365 ;
        RECT 132.670 280.720 141.490 281.365 ;
        RECT 142.330 280.720 151.150 281.365 ;
        RECT 151.990 280.720 160.810 281.365 ;
        RECT 161.650 280.720 170.470 281.365 ;
        RECT 171.310 280.720 180.130 281.365 ;
        RECT 180.970 280.720 189.790 281.365 ;
        RECT 190.630 280.720 199.450 281.365 ;
        RECT 200.290 280.720 209.110 281.365 ;
        RECT 209.950 280.720 218.770 281.365 ;
        RECT 219.610 280.720 228.430 281.365 ;
        RECT 229.270 280.720 238.090 281.365 ;
        RECT 238.930 280.720 247.750 281.365 ;
        RECT 3.320 4.280 248.310 280.720 ;
        RECT 3.870 3.555 6.250 4.280 ;
        RECT 7.090 3.555 9.470 4.280 ;
        RECT 10.310 3.555 12.690 4.280 ;
        RECT 13.530 3.555 15.910 4.280 ;
        RECT 16.750 3.555 19.130 4.280 ;
        RECT 19.970 3.555 22.350 4.280 ;
        RECT 23.190 3.555 25.570 4.280 ;
        RECT 26.410 3.555 28.790 4.280 ;
        RECT 29.630 3.555 32.010 4.280 ;
        RECT 32.850 3.555 35.230 4.280 ;
        RECT 36.070 3.555 38.450 4.280 ;
        RECT 39.290 3.555 41.670 4.280 ;
        RECT 42.510 3.555 44.890 4.280 ;
        RECT 45.730 3.555 48.110 4.280 ;
        RECT 48.950 3.555 51.330 4.280 ;
        RECT 52.170 3.555 54.550 4.280 ;
        RECT 55.390 3.555 57.770 4.280 ;
        RECT 58.610 3.555 60.990 4.280 ;
        RECT 61.830 3.555 64.210 4.280 ;
        RECT 65.050 3.555 67.430 4.280 ;
        RECT 68.270 3.555 70.650 4.280 ;
        RECT 71.490 3.555 73.870 4.280 ;
        RECT 74.710 3.555 77.090 4.280 ;
        RECT 77.930 3.555 80.310 4.280 ;
        RECT 81.150 3.555 83.530 4.280 ;
        RECT 84.370 3.555 86.750 4.280 ;
        RECT 87.590 3.555 89.970 4.280 ;
        RECT 90.810 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.410 4.280 ;
        RECT 97.250 3.555 99.630 4.280 ;
        RECT 100.470 3.555 102.850 4.280 ;
        RECT 103.690 3.555 106.070 4.280 ;
        RECT 106.910 3.555 109.290 4.280 ;
        RECT 110.130 3.555 112.510 4.280 ;
        RECT 113.350 3.555 115.730 4.280 ;
        RECT 116.570 3.555 118.950 4.280 ;
        RECT 119.790 3.555 122.170 4.280 ;
        RECT 123.010 3.555 125.390 4.280 ;
        RECT 126.230 3.555 128.610 4.280 ;
        RECT 129.450 3.555 131.830 4.280 ;
        RECT 132.670 3.555 135.050 4.280 ;
        RECT 135.890 3.555 138.270 4.280 ;
        RECT 139.110 3.555 141.490 4.280 ;
        RECT 142.330 3.555 144.710 4.280 ;
        RECT 145.550 3.555 147.930 4.280 ;
        RECT 148.770 3.555 151.150 4.280 ;
        RECT 151.990 3.555 154.370 4.280 ;
        RECT 155.210 3.555 157.590 4.280 ;
        RECT 158.430 3.555 160.810 4.280 ;
        RECT 161.650 3.555 164.030 4.280 ;
        RECT 164.870 3.555 167.250 4.280 ;
        RECT 168.090 3.555 170.470 4.280 ;
        RECT 171.310 3.555 173.690 4.280 ;
        RECT 174.530 3.555 176.910 4.280 ;
        RECT 177.750 3.555 180.130 4.280 ;
        RECT 180.970 3.555 183.350 4.280 ;
        RECT 184.190 3.555 186.570 4.280 ;
        RECT 187.410 3.555 189.790 4.280 ;
        RECT 190.630 3.555 193.010 4.280 ;
        RECT 193.850 3.555 196.230 4.280 ;
        RECT 197.070 3.555 199.450 4.280 ;
        RECT 200.290 3.555 202.670 4.280 ;
        RECT 203.510 3.555 205.890 4.280 ;
        RECT 206.730 3.555 209.110 4.280 ;
        RECT 209.950 3.555 212.330 4.280 ;
        RECT 213.170 3.555 215.550 4.280 ;
        RECT 216.390 3.555 218.770 4.280 ;
        RECT 219.610 3.555 221.990 4.280 ;
        RECT 222.830 3.555 225.210 4.280 ;
        RECT 226.050 3.555 228.430 4.280 ;
        RECT 229.270 3.555 231.650 4.280 ;
        RECT 232.490 3.555 234.870 4.280 ;
        RECT 235.710 3.555 238.090 4.280 ;
        RECT 238.930 3.555 241.310 4.280 ;
        RECT 242.150 3.555 244.530 4.280 ;
        RECT 245.370 3.555 247.750 4.280 ;
      LAYER met3 ;
        RECT 4.000 280.480 250.600 281.345 ;
        RECT 4.000 279.840 251.000 280.480 ;
        RECT 4.400 278.440 251.000 279.840 ;
        RECT 4.000 277.800 251.000 278.440 ;
        RECT 4.000 276.400 250.600 277.800 ;
        RECT 4.000 275.760 251.000 276.400 ;
        RECT 4.400 274.360 251.000 275.760 ;
        RECT 4.000 273.720 251.000 274.360 ;
        RECT 4.000 272.320 250.600 273.720 ;
        RECT 4.000 271.680 251.000 272.320 ;
        RECT 4.400 270.280 251.000 271.680 ;
        RECT 4.000 269.640 251.000 270.280 ;
        RECT 4.000 268.240 250.600 269.640 ;
        RECT 4.000 267.600 251.000 268.240 ;
        RECT 4.400 266.200 251.000 267.600 ;
        RECT 4.000 265.560 251.000 266.200 ;
        RECT 4.000 264.160 250.600 265.560 ;
        RECT 4.000 263.520 251.000 264.160 ;
        RECT 4.400 262.120 251.000 263.520 ;
        RECT 4.000 261.480 251.000 262.120 ;
        RECT 4.000 260.080 250.600 261.480 ;
        RECT 4.000 259.440 251.000 260.080 ;
        RECT 4.400 258.040 251.000 259.440 ;
        RECT 4.000 257.400 251.000 258.040 ;
        RECT 4.000 256.000 250.600 257.400 ;
        RECT 4.000 255.360 251.000 256.000 ;
        RECT 4.400 253.960 251.000 255.360 ;
        RECT 4.000 253.320 251.000 253.960 ;
        RECT 4.000 251.920 250.600 253.320 ;
        RECT 4.000 251.280 251.000 251.920 ;
        RECT 4.400 249.880 251.000 251.280 ;
        RECT 4.000 249.240 251.000 249.880 ;
        RECT 4.000 247.840 250.600 249.240 ;
        RECT 4.000 247.200 251.000 247.840 ;
        RECT 4.400 245.800 251.000 247.200 ;
        RECT 4.000 245.160 251.000 245.800 ;
        RECT 4.000 243.760 250.600 245.160 ;
        RECT 4.000 243.120 251.000 243.760 ;
        RECT 4.400 241.720 251.000 243.120 ;
        RECT 4.000 241.080 251.000 241.720 ;
        RECT 4.000 239.680 250.600 241.080 ;
        RECT 4.000 239.040 251.000 239.680 ;
        RECT 4.400 237.640 251.000 239.040 ;
        RECT 4.000 237.000 251.000 237.640 ;
        RECT 4.000 235.600 250.600 237.000 ;
        RECT 4.000 234.960 251.000 235.600 ;
        RECT 4.400 233.560 251.000 234.960 ;
        RECT 4.000 232.920 251.000 233.560 ;
        RECT 4.000 231.520 250.600 232.920 ;
        RECT 4.000 230.880 251.000 231.520 ;
        RECT 4.400 229.480 251.000 230.880 ;
        RECT 4.000 228.840 251.000 229.480 ;
        RECT 4.000 227.440 250.600 228.840 ;
        RECT 4.000 226.800 251.000 227.440 ;
        RECT 4.400 225.400 251.000 226.800 ;
        RECT 4.000 224.760 251.000 225.400 ;
        RECT 4.000 223.360 250.600 224.760 ;
        RECT 4.000 222.720 251.000 223.360 ;
        RECT 4.400 221.320 251.000 222.720 ;
        RECT 4.000 220.680 251.000 221.320 ;
        RECT 4.000 219.280 250.600 220.680 ;
        RECT 4.000 218.640 251.000 219.280 ;
        RECT 4.400 217.240 251.000 218.640 ;
        RECT 4.000 216.600 251.000 217.240 ;
        RECT 4.000 215.200 250.600 216.600 ;
        RECT 4.000 214.560 251.000 215.200 ;
        RECT 4.400 213.160 251.000 214.560 ;
        RECT 4.000 212.520 251.000 213.160 ;
        RECT 4.000 211.120 250.600 212.520 ;
        RECT 4.000 210.480 251.000 211.120 ;
        RECT 4.400 209.080 251.000 210.480 ;
        RECT 4.000 208.440 251.000 209.080 ;
        RECT 4.000 207.040 250.600 208.440 ;
        RECT 4.000 206.400 251.000 207.040 ;
        RECT 4.400 205.000 251.000 206.400 ;
        RECT 4.000 204.360 251.000 205.000 ;
        RECT 4.000 202.960 250.600 204.360 ;
        RECT 4.000 202.320 251.000 202.960 ;
        RECT 4.400 200.920 251.000 202.320 ;
        RECT 4.000 200.280 251.000 200.920 ;
        RECT 4.000 198.880 250.600 200.280 ;
        RECT 4.000 198.240 251.000 198.880 ;
        RECT 4.400 196.840 251.000 198.240 ;
        RECT 4.000 196.200 251.000 196.840 ;
        RECT 4.000 194.800 250.600 196.200 ;
        RECT 4.000 194.160 251.000 194.800 ;
        RECT 4.400 192.760 251.000 194.160 ;
        RECT 4.000 192.120 251.000 192.760 ;
        RECT 4.000 190.720 250.600 192.120 ;
        RECT 4.000 190.080 251.000 190.720 ;
        RECT 4.400 188.680 251.000 190.080 ;
        RECT 4.000 188.040 251.000 188.680 ;
        RECT 4.000 186.640 250.600 188.040 ;
        RECT 4.000 186.000 251.000 186.640 ;
        RECT 4.400 184.600 251.000 186.000 ;
        RECT 4.000 183.960 251.000 184.600 ;
        RECT 4.000 182.560 250.600 183.960 ;
        RECT 4.000 181.920 251.000 182.560 ;
        RECT 4.400 180.520 251.000 181.920 ;
        RECT 4.000 179.880 251.000 180.520 ;
        RECT 4.000 178.480 250.600 179.880 ;
        RECT 4.000 177.840 251.000 178.480 ;
        RECT 4.400 176.440 251.000 177.840 ;
        RECT 4.000 175.800 251.000 176.440 ;
        RECT 4.000 174.400 250.600 175.800 ;
        RECT 4.000 173.760 251.000 174.400 ;
        RECT 4.400 172.360 251.000 173.760 ;
        RECT 4.000 171.720 251.000 172.360 ;
        RECT 4.000 170.320 250.600 171.720 ;
        RECT 4.000 169.680 251.000 170.320 ;
        RECT 4.400 168.280 251.000 169.680 ;
        RECT 4.000 167.640 251.000 168.280 ;
        RECT 4.000 166.240 250.600 167.640 ;
        RECT 4.000 165.600 251.000 166.240 ;
        RECT 4.400 164.200 251.000 165.600 ;
        RECT 4.000 163.560 251.000 164.200 ;
        RECT 4.000 162.160 250.600 163.560 ;
        RECT 4.000 161.520 251.000 162.160 ;
        RECT 4.400 160.120 251.000 161.520 ;
        RECT 4.000 159.480 251.000 160.120 ;
        RECT 4.000 158.080 250.600 159.480 ;
        RECT 4.000 157.440 251.000 158.080 ;
        RECT 4.400 156.040 251.000 157.440 ;
        RECT 4.000 155.400 251.000 156.040 ;
        RECT 4.000 154.000 250.600 155.400 ;
        RECT 4.000 153.360 251.000 154.000 ;
        RECT 4.400 151.960 251.000 153.360 ;
        RECT 4.000 151.320 251.000 151.960 ;
        RECT 4.000 149.920 250.600 151.320 ;
        RECT 4.000 149.280 251.000 149.920 ;
        RECT 4.400 147.880 251.000 149.280 ;
        RECT 4.000 147.240 251.000 147.880 ;
        RECT 4.000 145.840 250.600 147.240 ;
        RECT 4.000 145.200 251.000 145.840 ;
        RECT 4.400 143.800 251.000 145.200 ;
        RECT 4.000 143.160 251.000 143.800 ;
        RECT 4.000 141.760 250.600 143.160 ;
        RECT 4.000 141.120 251.000 141.760 ;
        RECT 4.400 139.720 251.000 141.120 ;
        RECT 4.000 139.080 251.000 139.720 ;
        RECT 4.000 137.680 250.600 139.080 ;
        RECT 4.000 137.040 251.000 137.680 ;
        RECT 4.400 135.640 251.000 137.040 ;
        RECT 4.000 135.000 251.000 135.640 ;
        RECT 4.000 133.600 250.600 135.000 ;
        RECT 4.000 132.960 251.000 133.600 ;
        RECT 4.400 131.560 251.000 132.960 ;
        RECT 4.000 130.920 251.000 131.560 ;
        RECT 4.000 129.520 250.600 130.920 ;
        RECT 4.000 128.880 251.000 129.520 ;
        RECT 4.400 127.480 251.000 128.880 ;
        RECT 4.000 126.840 251.000 127.480 ;
        RECT 4.000 125.440 250.600 126.840 ;
        RECT 4.000 124.800 251.000 125.440 ;
        RECT 4.400 123.400 251.000 124.800 ;
        RECT 4.000 122.760 251.000 123.400 ;
        RECT 4.000 121.360 250.600 122.760 ;
        RECT 4.000 120.720 251.000 121.360 ;
        RECT 4.400 119.320 251.000 120.720 ;
        RECT 4.000 118.680 251.000 119.320 ;
        RECT 4.000 117.280 250.600 118.680 ;
        RECT 4.000 116.640 251.000 117.280 ;
        RECT 4.400 115.240 251.000 116.640 ;
        RECT 4.000 114.600 251.000 115.240 ;
        RECT 4.000 113.200 250.600 114.600 ;
        RECT 4.000 112.560 251.000 113.200 ;
        RECT 4.400 111.160 251.000 112.560 ;
        RECT 4.000 110.520 251.000 111.160 ;
        RECT 4.000 109.120 250.600 110.520 ;
        RECT 4.000 108.480 251.000 109.120 ;
        RECT 4.400 107.080 251.000 108.480 ;
        RECT 4.000 106.440 251.000 107.080 ;
        RECT 4.000 105.040 250.600 106.440 ;
        RECT 4.000 104.400 251.000 105.040 ;
        RECT 4.400 103.000 251.000 104.400 ;
        RECT 4.000 102.360 251.000 103.000 ;
        RECT 4.000 100.960 250.600 102.360 ;
        RECT 4.000 100.320 251.000 100.960 ;
        RECT 4.400 98.920 251.000 100.320 ;
        RECT 4.000 98.280 251.000 98.920 ;
        RECT 4.000 96.880 250.600 98.280 ;
        RECT 4.000 96.240 251.000 96.880 ;
        RECT 4.400 94.840 251.000 96.240 ;
        RECT 4.000 94.200 251.000 94.840 ;
        RECT 4.000 92.800 250.600 94.200 ;
        RECT 4.000 92.160 251.000 92.800 ;
        RECT 4.400 90.760 251.000 92.160 ;
        RECT 4.000 90.120 251.000 90.760 ;
        RECT 4.000 88.720 250.600 90.120 ;
        RECT 4.000 88.080 251.000 88.720 ;
        RECT 4.400 86.680 251.000 88.080 ;
        RECT 4.000 86.040 251.000 86.680 ;
        RECT 4.000 84.640 250.600 86.040 ;
        RECT 4.000 84.000 251.000 84.640 ;
        RECT 4.400 82.600 251.000 84.000 ;
        RECT 4.000 81.960 251.000 82.600 ;
        RECT 4.000 80.560 250.600 81.960 ;
        RECT 4.000 79.920 251.000 80.560 ;
        RECT 4.400 78.520 251.000 79.920 ;
        RECT 4.000 77.880 251.000 78.520 ;
        RECT 4.000 76.480 250.600 77.880 ;
        RECT 4.000 75.840 251.000 76.480 ;
        RECT 4.400 74.440 251.000 75.840 ;
        RECT 4.000 73.800 251.000 74.440 ;
        RECT 4.000 72.400 250.600 73.800 ;
        RECT 4.000 71.760 251.000 72.400 ;
        RECT 4.400 70.360 251.000 71.760 ;
        RECT 4.000 69.720 251.000 70.360 ;
        RECT 4.000 68.320 250.600 69.720 ;
        RECT 4.000 67.680 251.000 68.320 ;
        RECT 4.400 66.280 251.000 67.680 ;
        RECT 4.000 65.640 251.000 66.280 ;
        RECT 4.000 64.240 250.600 65.640 ;
        RECT 4.000 63.600 251.000 64.240 ;
        RECT 4.400 62.200 251.000 63.600 ;
        RECT 4.000 61.560 251.000 62.200 ;
        RECT 4.000 60.160 250.600 61.560 ;
        RECT 4.000 59.520 251.000 60.160 ;
        RECT 4.400 58.120 251.000 59.520 ;
        RECT 4.000 57.480 251.000 58.120 ;
        RECT 4.000 56.080 250.600 57.480 ;
        RECT 4.000 55.440 251.000 56.080 ;
        RECT 4.400 54.040 251.000 55.440 ;
        RECT 4.000 53.400 251.000 54.040 ;
        RECT 4.000 52.000 250.600 53.400 ;
        RECT 4.000 51.360 251.000 52.000 ;
        RECT 4.400 49.960 251.000 51.360 ;
        RECT 4.000 49.320 251.000 49.960 ;
        RECT 4.000 47.920 250.600 49.320 ;
        RECT 4.000 47.280 251.000 47.920 ;
        RECT 4.400 45.880 251.000 47.280 ;
        RECT 4.000 45.240 251.000 45.880 ;
        RECT 4.000 43.840 250.600 45.240 ;
        RECT 4.000 43.200 251.000 43.840 ;
        RECT 4.400 41.800 251.000 43.200 ;
        RECT 4.000 41.160 251.000 41.800 ;
        RECT 4.000 39.760 250.600 41.160 ;
        RECT 4.000 39.120 251.000 39.760 ;
        RECT 4.400 37.720 251.000 39.120 ;
        RECT 4.000 37.080 251.000 37.720 ;
        RECT 4.000 35.680 250.600 37.080 ;
        RECT 4.000 35.040 251.000 35.680 ;
        RECT 4.400 33.640 251.000 35.040 ;
        RECT 4.000 33.000 251.000 33.640 ;
        RECT 4.000 31.600 250.600 33.000 ;
        RECT 4.000 30.960 251.000 31.600 ;
        RECT 4.400 29.560 251.000 30.960 ;
        RECT 4.000 28.920 251.000 29.560 ;
        RECT 4.000 27.520 250.600 28.920 ;
        RECT 4.000 26.880 251.000 27.520 ;
        RECT 4.400 25.480 251.000 26.880 ;
        RECT 4.000 24.840 251.000 25.480 ;
        RECT 4.000 23.440 250.600 24.840 ;
        RECT 4.000 22.800 251.000 23.440 ;
        RECT 4.400 21.400 251.000 22.800 ;
        RECT 4.000 20.760 251.000 21.400 ;
        RECT 4.000 19.360 250.600 20.760 ;
        RECT 4.000 18.720 251.000 19.360 ;
        RECT 4.400 17.320 251.000 18.720 ;
        RECT 4.000 16.680 251.000 17.320 ;
        RECT 4.000 15.280 250.600 16.680 ;
        RECT 4.000 14.640 251.000 15.280 ;
        RECT 4.400 13.240 251.000 14.640 ;
        RECT 4.000 12.600 251.000 13.240 ;
        RECT 4.000 11.200 250.600 12.600 ;
        RECT 4.000 10.560 251.000 11.200 ;
        RECT 4.400 9.160 251.000 10.560 ;
        RECT 4.000 8.520 251.000 9.160 ;
        RECT 4.000 7.120 250.600 8.520 ;
        RECT 4.000 6.480 251.000 7.120 ;
        RECT 4.400 5.080 251.000 6.480 ;
        RECT 4.000 4.440 251.000 5.080 ;
        RECT 4.000 3.575 250.600 4.440 ;
      LAYER met4 ;
        RECT 30.655 10.240 39.320 259.585 ;
        RECT 41.720 10.240 64.320 259.585 ;
        RECT 66.720 10.240 89.320 259.585 ;
        RECT 91.720 10.240 114.320 259.585 ;
        RECT 116.720 10.240 139.320 259.585 ;
        RECT 141.720 10.240 164.320 259.585 ;
        RECT 166.720 10.240 189.320 259.585 ;
        RECT 191.720 10.240 214.320 259.585 ;
        RECT 216.720 10.240 234.305 259.585 ;
        RECT 30.655 7.655 234.305 10.240 ;
  END
END top_tile
END LIBRARY

