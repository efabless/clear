magic
tech sky130A
magscale 1 2
timestamp 1682507126
<< viali >>
rect 3985 24361 4019 24395
rect 4169 24361 4203 24395
rect 4353 24361 4387 24395
rect 9137 24361 9171 24395
rect 24593 24361 24627 24395
rect 32965 24361 32999 24395
rect 38025 24361 38059 24395
rect 39313 24361 39347 24395
rect 40049 24361 40083 24395
rect 44741 24361 44775 24395
rect 1593 24293 1627 24327
rect 14289 24293 14323 24327
rect 18981 24293 19015 24327
rect 28917 24293 28951 24327
rect 46857 24293 46891 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 16865 24225 16899 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25237 24225 25271 24259
rect 26341 24225 26375 24259
rect 28365 24225 28399 24259
rect 29745 24225 29779 24259
rect 35541 24225 35575 24259
rect 38669 24225 38703 24259
rect 1777 24157 1811 24191
rect 2145 24157 2179 24191
rect 4629 24157 4663 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 14933 24157 14967 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 24961 24157 24995 24191
rect 26249 24157 26283 24191
rect 29101 24157 29135 24191
rect 30021 24157 30055 24191
rect 31033 24157 31067 24191
rect 32321 24157 32355 24191
rect 33425 24157 33459 24191
rect 34345 24157 34379 24191
rect 34897 24157 34931 24191
rect 36921 24157 36955 24191
rect 38485 24157 38519 24191
rect 39221 24157 39255 24191
rect 40233 24157 40267 24191
rect 41245 24157 41279 24191
rect 41521 24157 41555 24191
rect 42625 24157 42659 24191
rect 45201 24157 45235 24191
rect 45937 24157 45971 24191
rect 46673 24157 46707 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48513 24157 48547 24191
rect 49065 24157 49099 24191
rect 16129 24089 16163 24123
rect 17141 24089 17175 24123
rect 27353 24089 27387 24123
rect 36093 24089 36127 24123
rect 37565 24089 37599 24123
rect 40509 24089 40543 24123
rect 6561 24021 6595 24055
rect 11713 24021 11747 24055
rect 11805 24021 11839 24055
rect 11989 24021 12023 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 23857 24021 23891 24055
rect 25053 24021 25087 24055
rect 25789 24021 25823 24055
rect 26157 24021 26191 24055
rect 26985 24021 27019 24055
rect 27261 24021 27295 24055
rect 27721 24021 27755 24055
rect 28089 24021 28123 24055
rect 28181 24021 28215 24055
rect 31677 24021 31711 24055
rect 34069 24021 34103 24055
rect 36185 24021 36219 24055
rect 36737 24021 36771 24055
rect 37657 24021 37691 24055
rect 40693 24021 40727 24055
rect 40877 24021 40911 24055
rect 43913 24021 43947 24055
rect 45385 24021 45419 24055
rect 46121 24021 46155 24055
rect 47961 24021 47995 24055
rect 48697 24021 48731 24055
rect 16773 23817 16807 23851
rect 33977 23817 34011 23851
rect 36553 23817 36587 23851
rect 36921 23817 36955 23851
rect 37473 23817 37507 23851
rect 38945 23817 38979 23851
rect 42165 23817 42199 23851
rect 42441 23817 42475 23851
rect 42993 23817 43027 23851
rect 43269 23817 43303 23851
rect 45753 23817 45787 23851
rect 47593 23817 47627 23851
rect 7113 23749 7147 23783
rect 9137 23749 9171 23783
rect 10977 23749 11011 23783
rect 14289 23749 14323 23783
rect 18245 23749 18279 23783
rect 19165 23749 19199 23783
rect 21373 23749 21407 23783
rect 25145 23749 25179 23783
rect 30757 23749 30791 23783
rect 42809 23749 42843 23783
rect 43637 23749 43671 23783
rect 1685 23681 1719 23715
rect 2789 23681 2823 23715
rect 3985 23681 4019 23715
rect 4629 23681 4663 23715
rect 7205 23681 7239 23715
rect 8125 23681 8159 23715
rect 9873 23681 9907 23715
rect 11713 23681 11747 23715
rect 13277 23681 13311 23715
rect 15025 23681 15059 23715
rect 17233 23681 17267 23715
rect 21189 23681 21223 23715
rect 29653 23681 29687 23715
rect 30941 23681 30975 23715
rect 31585 23681 31619 23715
rect 32332 23681 32366 23715
rect 34621 23681 34655 23715
rect 35708 23681 35742 23715
rect 35909 23681 35943 23715
rect 36461 23681 36495 23715
rect 38301 23681 38335 23715
rect 38853 23681 38887 23715
rect 40049 23681 40083 23715
rect 40233 23681 40267 23715
rect 42625 23681 42659 23715
rect 44281 23681 44315 23715
rect 44833 23681 44867 23715
rect 46765 23681 46799 23715
rect 47317 23681 47351 23715
rect 48881 23681 48915 23715
rect 49157 23681 49191 23715
rect 5457 23613 5491 23647
rect 7389 23613 7423 23647
rect 11989 23613 12023 23647
rect 16129 23613 16163 23647
rect 18889 23613 18923 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 24225 23613 24259 23647
rect 24869 23613 24903 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 29377 23613 29411 23647
rect 32965 23613 32999 23647
rect 34345 23613 34379 23647
rect 39497 23613 39531 23647
rect 40693 23613 40727 23647
rect 40969 23613 41003 23647
rect 41981 23613 42015 23647
rect 2329 23545 2363 23579
rect 26617 23545 26651 23579
rect 33425 23545 33459 23579
rect 33701 23545 33735 23579
rect 38117 23545 38151 23579
rect 41797 23545 41831 23579
rect 44465 23545 44499 23579
rect 6377 23477 6411 23511
rect 6745 23477 6779 23511
rect 20637 23477 20671 23511
rect 23765 23477 23799 23511
rect 28917 23477 28951 23511
rect 31401 23477 31435 23511
rect 31861 23477 31895 23511
rect 33241 23477 33275 23511
rect 33793 23477 33827 23511
rect 39313 23477 39347 23511
rect 43729 23477 43763 23511
rect 46949 23477 46983 23511
rect 48697 23477 48731 23511
rect 14473 23273 14507 23307
rect 25789 23273 25823 23307
rect 29009 23273 29043 23307
rect 34897 23273 34931 23307
rect 3433 23205 3467 23239
rect 9137 23205 9171 23239
rect 11161 23205 11195 23239
rect 18889 23205 18923 23239
rect 21833 23205 21867 23239
rect 24685 23205 24719 23239
rect 34161 23205 34195 23239
rect 36829 23205 36863 23239
rect 40693 23205 40727 23239
rect 3617 23137 3651 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 11713 23137 11747 23171
rect 20085 23137 20119 23171
rect 22293 23137 22327 23171
rect 25237 23137 25271 23171
rect 26433 23137 26467 23171
rect 27261 23137 27295 23171
rect 29285 23137 29319 23171
rect 29745 23137 29779 23171
rect 30021 23137 30055 23171
rect 39497 23137 39531 23171
rect 42441 23137 42475 23171
rect 1777 23069 1811 23103
rect 3985 23069 4019 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9413 23069 9447 23103
rect 14381 23069 14415 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 26249 23069 26283 23103
rect 31953 23069 31987 23103
rect 33057 23069 33091 23103
rect 34345 23069 34379 23103
rect 35081 23069 35115 23103
rect 35541 23069 35575 23103
rect 35817 23069 35851 23103
rect 37013 23069 37047 23103
rect 38485 23069 38519 23103
rect 38945 23069 38979 23103
rect 40233 23069 40267 23103
rect 40877 23069 40911 23103
rect 41521 23069 41555 23103
rect 42165 23069 42199 23103
rect 2789 23001 2823 23035
rect 9689 23001 9723 23035
rect 11989 23001 12023 23035
rect 13829 23001 13863 23035
rect 16497 23001 16531 23035
rect 17417 23001 17451 23035
rect 20361 23001 20395 23035
rect 22569 23001 22603 23035
rect 24961 23001 24995 23035
rect 26801 23001 26835 23035
rect 27537 23001 27571 23035
rect 37565 23001 37599 23035
rect 38301 23001 38335 23035
rect 4215 22933 4249 22967
rect 13461 22933 13495 22967
rect 14933 22933 14967 22967
rect 19441 22933 19475 22967
rect 24041 22933 24075 22967
rect 25145 22933 25179 22967
rect 26157 22933 26191 22967
rect 31493 22933 31527 22967
rect 32597 22933 32631 22967
rect 33701 22933 33735 22967
rect 37657 22933 37691 22967
rect 39129 22933 39163 22967
rect 40049 22933 40083 22967
rect 41337 22933 41371 22967
rect 41981 22933 42015 22967
rect 18613 22729 18647 22763
rect 19073 22729 19107 22763
rect 24869 22729 24903 22763
rect 25697 22729 25731 22763
rect 26801 22729 26835 22763
rect 31585 22729 31619 22763
rect 32965 22729 32999 22763
rect 33333 22729 33367 22763
rect 37473 22729 37507 22763
rect 39957 22729 39991 22763
rect 40141 22729 40175 22763
rect 41153 22729 41187 22763
rect 5549 22661 5583 22695
rect 6653 22661 6687 22695
rect 7113 22661 7147 22695
rect 10701 22661 10735 22695
rect 11805 22661 11839 22695
rect 12725 22661 12759 22695
rect 16129 22661 16163 22695
rect 16773 22661 16807 22695
rect 17141 22661 17175 22695
rect 19993 22661 20027 22695
rect 23397 22661 23431 22695
rect 37289 22661 37323 22695
rect 40417 22661 40451 22695
rect 1777 22593 1811 22627
rect 3525 22593 3559 22627
rect 4629 22593 4663 22627
rect 7205 22593 7239 22627
rect 7941 22593 7975 22627
rect 9781 22593 9815 22627
rect 12449 22593 12483 22627
rect 14933 22593 14967 22627
rect 19717 22593 19751 22627
rect 22017 22593 22051 22627
rect 23121 22593 23155 22627
rect 27169 22593 27203 22627
rect 28365 22593 28399 22627
rect 30941 22593 30975 22627
rect 31861 22593 31895 22627
rect 32321 22593 32355 22627
rect 33885 22593 33919 22627
rect 34621 22593 34655 22627
rect 35725 22593 35759 22627
rect 36461 22593 36495 22627
rect 2789 22525 2823 22559
rect 4169 22525 4203 22559
rect 7389 22525 7423 22559
rect 8677 22525 8711 22559
rect 16865 22525 16899 22559
rect 25789 22525 25823 22559
rect 25881 22525 25915 22559
rect 28641 22525 28675 22559
rect 31033 22525 31067 22559
rect 31125 22525 31159 22559
rect 34345 22525 34379 22559
rect 35909 22525 35943 22559
rect 37933 22525 37967 22559
rect 38209 22525 38243 22559
rect 6745 22457 6779 22491
rect 11989 22457 12023 22491
rect 26341 22457 26375 22491
rect 30573 22457 30607 22491
rect 33701 22457 33735 22491
rect 40509 22457 40543 22491
rect 6469 22389 6503 22423
rect 14197 22389 14231 22423
rect 14565 22389 14599 22423
rect 21465 22389 21499 22423
rect 22661 22389 22695 22423
rect 25329 22389 25363 22423
rect 26617 22389 26651 22423
rect 27813 22389 27847 22423
rect 30113 22389 30147 22423
rect 36553 22389 36587 22423
rect 36921 22389 36955 22423
rect 39681 22389 39715 22423
rect 17404 22185 17438 22219
rect 20085 22185 20119 22219
rect 26052 22185 26086 22219
rect 29285 22185 29319 22219
rect 29561 22185 29595 22219
rect 37565 22185 37599 22219
rect 14105 22117 14139 22151
rect 23305 22117 23339 22151
rect 27537 22117 27571 22151
rect 34345 22117 34379 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 7297 22049 7331 22083
rect 8769 22049 8803 22083
rect 9781 22049 9815 22083
rect 9965 22049 9999 22083
rect 11253 22049 11287 22083
rect 13369 22049 13403 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20821 22049 20855 22083
rect 23949 22049 23983 22083
rect 25237 22049 25271 22083
rect 30481 22049 30515 22083
rect 30665 22049 30699 22083
rect 32965 22049 32999 22083
rect 35173 22049 35207 22083
rect 39681 22049 39715 22083
rect 1777 21981 1811 22015
rect 4077 21981 4111 22015
rect 6377 21981 6411 22015
rect 6837 21981 6871 22015
rect 10609 21981 10643 22015
rect 12357 21981 12391 22015
rect 14565 21981 14599 22015
rect 15393 21981 15427 22015
rect 20361 21981 20395 22015
rect 22201 21981 22235 22015
rect 23673 21981 23707 22015
rect 23765 21981 23799 22015
rect 25789 21981 25823 22015
rect 27997 21981 28031 22015
rect 31217 21981 31251 22015
rect 32321 21981 32355 22015
rect 33425 21981 33459 22015
rect 37105 21981 37139 22015
rect 37749 21981 37783 22015
rect 38393 21981 38427 22015
rect 39037 21981 39071 22015
rect 39313 21981 39347 22015
rect 5641 21913 5675 21947
rect 9045 21913 9079 21947
rect 19533 21913 19567 21947
rect 25053 21913 25087 21947
rect 34989 21913 35023 21947
rect 35725 21913 35759 21947
rect 35909 21913 35943 21947
rect 36921 21913 36955 21947
rect 3433 21845 3467 21879
rect 3617 21845 3651 21879
rect 5917 21845 5951 21879
rect 6193 21845 6227 21879
rect 8493 21845 8527 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 14657 21845 14691 21879
rect 18889 21845 18923 21879
rect 19625 21845 19659 21879
rect 22845 21845 22879 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 28641 21845 28675 21879
rect 29009 21845 29043 21879
rect 29101 21845 29135 21879
rect 30021 21845 30055 21879
rect 30389 21845 30423 21879
rect 31861 21845 31895 21879
rect 34069 21845 34103 21879
rect 36185 21845 36219 21879
rect 36369 21845 36403 21879
rect 38209 21845 38243 21879
rect 38853 21845 38887 21879
rect 7113 21641 7147 21675
rect 9597 21641 9631 21675
rect 10149 21641 10183 21675
rect 11989 21641 12023 21675
rect 15945 21641 15979 21675
rect 17785 21641 17819 21675
rect 22477 21641 22511 21675
rect 25973 21641 26007 21675
rect 27261 21641 27295 21675
rect 27721 21641 27755 21675
rect 30665 21641 30699 21675
rect 31033 21641 31067 21675
rect 31125 21641 31159 21675
rect 33425 21641 33459 21675
rect 34713 21641 34747 21675
rect 35909 21641 35943 21675
rect 36001 21641 36035 21675
rect 37473 21641 37507 21675
rect 38393 21641 38427 21675
rect 5733 21573 5767 21607
rect 8125 21573 8159 21607
rect 23673 21573 23707 21607
rect 26065 21573 26099 21607
rect 34069 21573 34103 21607
rect 37289 21573 37323 21607
rect 38301 21573 38335 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 5641 21505 5675 21539
rect 7021 21505 7055 21539
rect 7481 21505 7515 21539
rect 10793 21505 10827 21539
rect 12357 21505 12391 21539
rect 13185 21505 13219 21539
rect 15209 21505 15243 21539
rect 16681 21505 16715 21539
rect 20821 21505 20855 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 27629 21505 27663 21539
rect 31769 21505 31803 21539
rect 32321 21505 32355 21539
rect 34621 21505 34655 21539
rect 35357 21505 35391 21539
rect 36829 21505 36863 21539
rect 37841 21505 37875 21539
rect 47961 21505 47995 21539
rect 2789 21437 2823 21471
rect 3893 21437 3927 21471
rect 5917 21437 5951 21471
rect 7205 21437 7239 21471
rect 7849 21437 7883 21471
rect 10885 21437 10919 21471
rect 10977 21437 11011 21471
rect 12449 21437 12483 21471
rect 12541 21437 12575 21471
rect 13461 21437 13495 21471
rect 14933 21437 14967 21471
rect 16037 21437 16071 21471
rect 16129 21437 16163 21471
rect 16957 21437 16991 21471
rect 17877 21437 17911 21471
rect 17969 21437 18003 21471
rect 18613 21437 18647 21471
rect 18889 21437 18923 21471
rect 22661 21437 22695 21471
rect 25145 21437 25179 21471
rect 26157 21437 26191 21471
rect 27813 21437 27847 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 33885 21437 33919 21471
rect 35541 21437 35575 21471
rect 49157 21437 49191 21471
rect 6653 21369 6687 21403
rect 26709 21369 26743 21403
rect 30205 21369 30239 21403
rect 31953 21369 31987 21403
rect 36645 21369 36679 21403
rect 37657 21369 37691 21403
rect 5273 21301 5307 21335
rect 6469 21301 6503 21335
rect 10425 21301 10459 21335
rect 11621 21301 11655 21335
rect 15577 21301 15611 21335
rect 17141 21301 17175 21335
rect 17417 21301 17451 21335
rect 20361 21301 20395 21335
rect 21465 21301 21499 21335
rect 22017 21301 22051 21335
rect 23121 21301 23155 21335
rect 25605 21301 25639 21335
rect 32965 21301 32999 21335
rect 38025 21301 38059 21335
rect 47593 21301 47627 21335
rect 5825 21097 5859 21131
rect 8033 21097 8067 21131
rect 19073 21097 19107 21131
rect 23029 21097 23063 21131
rect 27721 21097 27755 21131
rect 29285 21097 29319 21131
rect 31861 21097 31895 21131
rect 34161 21097 34195 21131
rect 37381 21097 37415 21131
rect 3433 21029 3467 21063
rect 8769 21029 8803 21063
rect 13737 21029 13771 21063
rect 35909 21029 35943 21063
rect 4445 20961 4479 20995
rect 6285 20961 6319 20995
rect 8309 20961 8343 20995
rect 12449 20961 12483 20995
rect 13829 20961 13863 20995
rect 14289 20961 14323 20995
rect 14473 20961 14507 20995
rect 15209 20961 15243 20995
rect 15393 20961 15427 20995
rect 16405 20961 16439 20995
rect 16497 20961 16531 20995
rect 17601 20961 17635 20995
rect 19441 20961 19475 20995
rect 22385 20961 22419 20995
rect 23489 20961 23523 20995
rect 23673 20961 23707 20995
rect 25145 20961 25179 20995
rect 25329 20961 25363 20995
rect 32229 20961 32263 20995
rect 32873 20961 32907 20995
rect 33149 20961 33183 20995
rect 1777 20893 1811 20927
rect 3985 20893 4019 20927
rect 9321 20893 9355 20927
rect 11621 20893 11655 20927
rect 12173 20893 12207 20927
rect 15117 20893 15151 20927
rect 16313 20893 16347 20927
rect 17141 20893 17175 20927
rect 25973 20893 26007 20927
rect 28181 20893 28215 20927
rect 29193 20893 29227 20927
rect 29745 20893 29779 20927
rect 30849 20893 30883 20927
rect 34345 20893 34379 20927
rect 2789 20825 2823 20859
rect 6561 20825 6595 20859
rect 10057 20825 10091 20859
rect 11069 20825 11103 20859
rect 19724 20825 19758 20859
rect 21649 20825 21683 20859
rect 23397 20825 23431 20859
rect 25053 20825 25087 20859
rect 26249 20825 26283 20859
rect 34989 20825 35023 20859
rect 35725 20825 35759 20859
rect 36461 20825 36495 20859
rect 36921 20825 36955 20859
rect 3617 20757 3651 20791
rect 5917 20757 5951 20791
rect 8493 20757 8527 20791
rect 11161 20757 11195 20791
rect 14749 20757 14783 20791
rect 15945 20757 15979 20791
rect 18797 20757 18831 20791
rect 21189 20757 21223 20791
rect 24225 20757 24259 20791
rect 24685 20757 24719 20791
rect 28825 20757 28859 20791
rect 30389 20757 30423 20791
rect 31493 20757 31527 20791
rect 35081 20757 35115 20791
rect 36553 20757 36587 20791
rect 37105 20757 37139 20791
rect 5641 20553 5675 20587
rect 11069 20553 11103 20587
rect 11989 20553 12023 20587
rect 13001 20553 13035 20587
rect 16681 20553 16715 20587
rect 17509 20553 17543 20587
rect 18153 20553 18187 20587
rect 18981 20553 19015 20587
rect 23581 20553 23615 20587
rect 27169 20553 27203 20587
rect 31769 20553 31803 20587
rect 31861 20553 31895 20587
rect 33241 20553 33275 20587
rect 35633 20553 35667 20587
rect 11897 20485 11931 20519
rect 12909 20485 12943 20519
rect 14013 20485 14047 20519
rect 23489 20485 23523 20519
rect 24593 20485 24627 20519
rect 26433 20485 26467 20519
rect 28733 20485 28767 20519
rect 34437 20485 34471 20519
rect 35081 20485 35115 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5733 20417 5767 20451
rect 6561 20417 6595 20451
rect 10977 20417 11011 20451
rect 13737 20417 13771 20451
rect 16037 20417 16071 20451
rect 17417 20417 17451 20451
rect 18889 20417 18923 20451
rect 19717 20417 19751 20451
rect 22017 20417 22051 20451
rect 26801 20417 26835 20451
rect 27537 20417 27571 20451
rect 28457 20417 28491 20451
rect 31033 20417 31067 20451
rect 31125 20417 31159 20451
rect 32321 20417 32355 20451
rect 33701 20417 33735 20451
rect 34897 20417 34931 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 5825 20349 5859 20383
rect 7021 20349 7055 20383
rect 8309 20349 8343 20383
rect 8585 20349 8619 20383
rect 8861 20349 8895 20383
rect 10333 20349 10367 20383
rect 13185 20349 13219 20383
rect 15485 20349 15519 20383
rect 17601 20349 17635 20383
rect 19165 20349 19199 20383
rect 21465 20349 21499 20383
rect 23765 20349 23799 20383
rect 24317 20349 24351 20383
rect 27629 20349 27663 20383
rect 27721 20349 27755 20383
rect 30205 20349 30239 20383
rect 31217 20349 31251 20383
rect 36001 20349 36035 20383
rect 16221 20281 16255 20315
rect 23121 20281 23155 20315
rect 26065 20281 26099 20315
rect 35909 20281 35943 20315
rect 5273 20213 5307 20247
rect 12541 20213 12575 20247
rect 17049 20213 17083 20247
rect 18521 20213 18555 20247
rect 19974 20213 20008 20247
rect 22661 20213 22695 20247
rect 26525 20213 26559 20247
rect 30665 20213 30699 20247
rect 32965 20213 32999 20247
rect 33793 20213 33827 20247
rect 34529 20213 34563 20247
rect 35265 20213 35299 20247
rect 35449 20213 35483 20247
rect 3617 20009 3651 20043
rect 4169 20009 4203 20043
rect 8953 20009 8987 20043
rect 17693 20009 17727 20043
rect 18153 20009 18187 20043
rect 21925 20009 21959 20043
rect 22385 20009 22419 20043
rect 26144 20009 26178 20043
rect 27629 20009 27663 20043
rect 34713 20009 34747 20043
rect 3893 19941 3927 19975
rect 14197 19941 14231 19975
rect 16405 19941 16439 19975
rect 3433 19873 3467 19907
rect 7573 19873 7607 19907
rect 10057 19873 10091 19907
rect 13645 19873 13679 19907
rect 14657 19873 14691 19907
rect 18705 19873 18739 19907
rect 19717 19873 19751 19907
rect 20177 19873 20211 19907
rect 20453 19873 20487 19907
rect 23673 19873 23707 19907
rect 25329 19873 25363 19907
rect 25881 19873 25915 19907
rect 29193 19873 29227 19907
rect 30021 19873 30055 19907
rect 31585 19873 31619 19907
rect 33517 19873 33551 19907
rect 33793 19873 33827 19907
rect 1777 19805 1811 19839
rect 4353 19805 4387 19839
rect 4905 19805 4939 19839
rect 7297 19805 7331 19839
rect 9413 19805 9447 19839
rect 17049 19805 17083 19839
rect 18613 19805 18647 19839
rect 22569 19805 22603 19839
rect 23397 19805 23431 19839
rect 23489 19805 23523 19839
rect 28089 19805 28123 19839
rect 29745 19805 29779 19839
rect 32229 19805 32263 19839
rect 33149 19805 33183 19839
rect 2789 19737 2823 19771
rect 5181 19737 5215 19771
rect 10333 19737 10367 19771
rect 12357 19737 12391 19771
rect 12541 19737 12575 19771
rect 14933 19737 14967 19771
rect 19533 19737 19567 19771
rect 25053 19737 25087 19771
rect 31401 19737 31435 19771
rect 31493 19737 31527 19771
rect 6653 19669 6687 19703
rect 9505 19669 9539 19703
rect 11805 19669 11839 19703
rect 13001 19669 13035 19703
rect 13369 19669 13403 19703
rect 13461 19669 13495 19703
rect 14381 19669 14415 19703
rect 18521 19669 18555 19703
rect 23029 19669 23063 19703
rect 24133 19669 24167 19703
rect 24685 19669 24719 19703
rect 25145 19669 25179 19703
rect 28733 19669 28767 19703
rect 29101 19669 29135 19703
rect 31033 19669 31067 19703
rect 32873 19669 32907 19703
rect 34897 19669 34931 19703
rect 3617 19465 3651 19499
rect 6009 19465 6043 19499
rect 9045 19465 9079 19499
rect 9781 19465 9815 19499
rect 10241 19465 10275 19499
rect 17877 19465 17911 19499
rect 18337 19465 18371 19499
rect 19073 19465 19107 19499
rect 21465 19465 21499 19499
rect 22477 19465 22511 19499
rect 22845 19465 22879 19499
rect 22937 19465 22971 19499
rect 24133 19465 24167 19499
rect 30113 19465 30147 19499
rect 14657 19397 14691 19431
rect 25789 19397 25823 19431
rect 31677 19397 31711 19431
rect 32413 19397 32447 19431
rect 33149 19397 33183 19431
rect 33609 19397 33643 19431
rect 1777 19329 1811 19363
rect 2789 19329 2823 19363
rect 3801 19329 3835 19363
rect 4261 19329 4295 19363
rect 6653 19329 6687 19363
rect 7297 19329 7331 19363
rect 9689 19329 9723 19363
rect 10149 19329 10183 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 13921 19329 13955 19363
rect 15669 19329 15703 19363
rect 15761 19329 15795 19363
rect 16957 19329 16991 19363
rect 18245 19329 18279 19363
rect 24041 19329 24075 19363
rect 24961 19329 24995 19363
rect 26617 19329 26651 19363
rect 27261 19329 27295 19363
rect 27905 19329 27939 19363
rect 28365 19329 28399 19363
rect 30573 19329 30607 19363
rect 31217 19329 31251 19363
rect 4537 19261 4571 19295
rect 7573 19261 7607 19295
rect 10425 19261 10459 19295
rect 11989 19261 12023 19295
rect 13461 19261 13495 19295
rect 15853 19261 15887 19295
rect 17509 19261 17543 19295
rect 18429 19261 18463 19295
rect 19717 19261 19751 19295
rect 19993 19261 20027 19295
rect 21925 19261 21959 19295
rect 23121 19261 23155 19295
rect 24225 19261 24259 19295
rect 28641 19261 28675 19295
rect 31585 19261 31619 19295
rect 31953 19261 31987 19295
rect 3341 19193 3375 19227
rect 6837 19193 6871 19227
rect 15301 19193 15335 19227
rect 23673 19193 23707 19227
rect 26433 19193 26467 19227
rect 9413 19125 9447 19159
rect 10977 19125 11011 19159
rect 16497 19125 16531 19159
rect 17049 19125 17083 19159
rect 22201 19125 22235 19159
rect 26249 19125 26283 19159
rect 32505 19125 32539 19159
rect 33241 19125 33275 19159
rect 3893 18921 3927 18955
rect 14289 18921 14323 18955
rect 18153 18921 18187 18955
rect 19349 18921 19383 18955
rect 25684 18921 25718 18955
rect 28825 18921 28859 18955
rect 32965 18921 32999 18955
rect 3617 18853 3651 18887
rect 4077 18853 4111 18887
rect 10609 18853 10643 18887
rect 11805 18853 11839 18887
rect 14565 18853 14599 18887
rect 17693 18853 17727 18887
rect 28641 18853 28675 18887
rect 32505 18853 32539 18887
rect 2053 18785 2087 18819
rect 3433 18785 3467 18819
rect 4997 18785 5031 18819
rect 5549 18785 5583 18819
rect 8401 18785 8435 18819
rect 9781 18785 9815 18819
rect 11253 18785 11287 18819
rect 12357 18785 12391 18819
rect 15209 18785 15243 18819
rect 18705 18785 18739 18819
rect 21189 18785 21223 18819
rect 21465 18785 21499 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 27169 18785 27203 18819
rect 28273 18785 28307 18819
rect 30297 18785 30331 18819
rect 1777 18717 1811 18751
rect 4721 18717 4755 18751
rect 7757 18717 7791 18751
rect 8217 18717 8251 18751
rect 9597 18717 9631 18751
rect 10977 18717 11011 18751
rect 13081 18717 13115 18751
rect 14749 18717 14783 18751
rect 18521 18717 18555 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 23397 18717 23431 18751
rect 29009 18717 29043 18751
rect 30205 18717 30239 18751
rect 30941 18717 30975 18751
rect 32689 18717 32723 18751
rect 5825 18649 5859 18683
rect 10517 18649 10551 18683
rect 11713 18649 11747 18683
rect 15485 18649 15519 18683
rect 17509 18649 17543 18683
rect 28089 18649 28123 18683
rect 30113 18649 30147 18683
rect 31953 18649 31987 18683
rect 4353 18581 4387 18615
rect 4813 18581 4847 18615
rect 7297 18581 7331 18615
rect 7849 18581 7883 18615
rect 8309 18581 8343 18615
rect 9229 18581 9263 18615
rect 9689 18581 9723 18615
rect 10333 18581 10367 18615
rect 11069 18581 11103 18615
rect 12173 18581 12207 18615
rect 12265 18581 12299 18615
rect 13737 18581 13771 18615
rect 16957 18581 16991 18615
rect 18613 18581 18647 18615
rect 20821 18581 20855 18615
rect 22937 18581 22971 18615
rect 24041 18581 24075 18615
rect 25053 18581 25087 18615
rect 27629 18581 27663 18615
rect 27997 18581 28031 18615
rect 29377 18581 29411 18615
rect 29745 18581 29779 18615
rect 31585 18581 31619 18615
rect 32137 18581 32171 18615
rect 5733 18377 5767 18411
rect 10149 18377 10183 18411
rect 10517 18377 10551 18411
rect 15669 18377 15703 18411
rect 15761 18377 15795 18411
rect 19809 18377 19843 18411
rect 27169 18377 27203 18411
rect 29837 18377 29871 18411
rect 30757 18377 30791 18411
rect 5641 18309 5675 18343
rect 11345 18309 11379 18343
rect 13921 18309 13955 18343
rect 17325 18309 17359 18343
rect 25329 18309 25363 18343
rect 31585 18309 31619 18343
rect 32137 18309 32171 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 8769 18241 8803 18275
rect 12081 18241 12115 18275
rect 13093 18241 13127 18275
rect 17233 18241 17267 18275
rect 18521 18241 18555 18275
rect 19533 18241 19567 18275
rect 20177 18241 20211 18275
rect 22017 18241 22051 18275
rect 23121 18241 23155 18275
rect 28089 18241 28123 18275
rect 30665 18241 30699 18275
rect 2053 18173 2087 18207
rect 3893 18173 3927 18207
rect 5917 18173 5951 18207
rect 6561 18173 6595 18207
rect 6837 18173 6871 18207
rect 9505 18173 9539 18207
rect 10609 18173 10643 18207
rect 10701 18173 10735 18207
rect 12265 18173 12299 18207
rect 13185 18173 13219 18207
rect 13277 18173 13311 18207
rect 14657 18173 14691 18207
rect 15945 18173 15979 18207
rect 17509 18173 17543 18207
rect 18613 18173 18647 18207
rect 18705 18173 18739 18207
rect 20269 18173 20303 18207
rect 20361 18173 20395 18207
rect 21281 18173 21315 18207
rect 22661 18173 22695 18207
rect 23397 18173 23431 18207
rect 26065 18173 26099 18207
rect 28365 18173 28399 18207
rect 30849 18173 30883 18207
rect 8309 18105 8343 18139
rect 12725 18105 12759 18139
rect 16865 18105 16899 18139
rect 24869 18105 24903 18139
rect 31769 18105 31803 18139
rect 5273 18037 5307 18071
rect 11621 18037 11655 18071
rect 15301 18037 15335 18071
rect 16405 18037 16439 18071
rect 18153 18037 18187 18071
rect 19349 18037 19383 18071
rect 21005 18037 21039 18071
rect 26709 18037 26743 18071
rect 27721 18037 27755 18071
rect 30297 18037 30331 18071
rect 3433 17833 3467 17867
rect 13921 17833 13955 17867
rect 14473 17833 14507 17867
rect 14841 17833 14875 17867
rect 18061 17833 18095 17867
rect 21741 17833 21775 17867
rect 21925 17833 21959 17867
rect 24685 17833 24719 17867
rect 26709 17833 26743 17867
rect 28917 17833 28951 17867
rect 31309 17833 31343 17867
rect 8769 17765 8803 17799
rect 2053 17697 2087 17731
rect 4445 17697 4479 17731
rect 6285 17697 6319 17731
rect 8217 17697 8251 17731
rect 10977 17697 11011 17731
rect 11069 17697 11103 17731
rect 11713 17697 11747 17731
rect 16313 17697 16347 17731
rect 16589 17697 16623 17731
rect 21189 17697 21223 17731
rect 21281 17697 21315 17731
rect 24409 17697 24443 17731
rect 24961 17697 24995 17731
rect 27169 17697 27203 17731
rect 30297 17697 30331 17731
rect 30849 17697 30883 17731
rect 1777 17629 1811 17663
rect 4077 17629 4111 17663
rect 6009 17629 6043 17663
rect 8033 17629 8067 17663
rect 15209 17629 15243 17663
rect 19349 17629 19383 17663
rect 19625 17629 19659 17663
rect 22293 17629 22327 17663
rect 29285 17629 29319 17663
rect 9137 17561 9171 17595
rect 9873 17561 9907 17595
rect 10425 17561 10459 17595
rect 11989 17561 12023 17595
rect 14381 17561 14415 17595
rect 18613 17561 18647 17595
rect 20269 17561 20303 17595
rect 22569 17561 22603 17595
rect 25237 17561 25271 17595
rect 27445 17561 27479 17595
rect 30113 17561 30147 17595
rect 31125 17561 31159 17595
rect 3617 17493 3651 17527
rect 7665 17493 7699 17527
rect 8125 17493 8159 17527
rect 10517 17493 10551 17527
rect 10885 17493 10919 17527
rect 13461 17493 13495 17527
rect 15853 17493 15887 17527
rect 18705 17493 18739 17527
rect 20729 17493 20763 17527
rect 21097 17493 21131 17527
rect 24041 17493 24075 17527
rect 29745 17493 29779 17527
rect 30205 17493 30239 17527
rect 30941 17493 30975 17527
rect 7205 17289 7239 17323
rect 7297 17289 7331 17323
rect 9597 17289 9631 17323
rect 9689 17289 9723 17323
rect 22569 17289 22603 17323
rect 22661 17289 22695 17323
rect 4353 17221 4387 17255
rect 11989 17221 12023 17255
rect 13737 17221 13771 17255
rect 18429 17221 18463 17255
rect 21833 17221 21867 17255
rect 23305 17221 23339 17255
rect 23949 17221 23983 17255
rect 24041 17221 24075 17255
rect 30021 17221 30055 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 5641 17153 5675 17187
rect 8401 17153 8435 17187
rect 10793 17153 10827 17187
rect 11805 17153 11839 17187
rect 12817 17153 12851 17187
rect 14749 17153 14783 17187
rect 14841 17153 14875 17187
rect 15669 17153 15703 17187
rect 17233 17153 17267 17187
rect 20177 17153 20211 17187
rect 20545 17153 20579 17187
rect 20821 17153 20855 17187
rect 24777 17153 24811 17187
rect 27905 17153 27939 17187
rect 2053 17085 2087 17119
rect 5733 17085 5767 17119
rect 5825 17085 5859 17119
rect 7389 17085 7423 17119
rect 8493 17085 8527 17119
rect 8677 17085 8711 17119
rect 9781 17085 9815 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 12909 17085 12943 17119
rect 13001 17085 13035 17119
rect 14933 17085 14967 17119
rect 17325 17085 17359 17119
rect 17509 17085 17543 17119
rect 18153 17085 18187 17119
rect 19901 17085 19935 17119
rect 22845 17085 22879 17119
rect 24133 17085 24167 17119
rect 25053 17085 25087 17119
rect 27261 17085 27295 17119
rect 28181 17085 28215 17119
rect 6837 17017 6871 17051
rect 12449 17017 12483 17051
rect 22201 17017 22235 17051
rect 5273 16949 5307 16983
rect 6469 16949 6503 16983
rect 8033 16949 8067 16983
rect 9229 16949 9263 16983
rect 10425 16949 10459 16983
rect 13829 16949 13863 16983
rect 14381 16949 14415 16983
rect 16313 16949 16347 16983
rect 16865 16949 16899 16983
rect 21465 16949 21499 16983
rect 23581 16949 23615 16983
rect 26525 16949 26559 16983
rect 29653 16949 29687 16983
rect 3433 16745 3467 16779
rect 10333 16745 10367 16779
rect 14473 16745 14507 16779
rect 16313 16745 16347 16779
rect 23305 16745 23339 16779
rect 3525 16677 3559 16711
rect 11805 16677 11839 16711
rect 13001 16677 13035 16711
rect 18797 16677 18831 16711
rect 6193 16609 6227 16643
rect 7113 16609 7147 16643
rect 7297 16609 7331 16643
rect 8309 16609 8343 16643
rect 8401 16609 8435 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 10241 16609 10275 16643
rect 12265 16609 12299 16643
rect 12449 16609 12483 16643
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 15669 16609 15703 16643
rect 19073 16609 19107 16643
rect 19441 16609 19475 16643
rect 22385 16609 22419 16643
rect 22477 16609 22511 16643
rect 23949 16609 23983 16643
rect 24501 16609 24535 16643
rect 25237 16609 25271 16643
rect 25421 16609 25455 16643
rect 25973 16609 26007 16643
rect 26249 16609 26283 16643
rect 27721 16609 27755 16643
rect 27813 16609 27847 16643
rect 28917 16609 28951 16643
rect 29101 16609 29135 16643
rect 30021 16609 30055 16643
rect 1777 16541 1811 16575
rect 4077 16541 4111 16575
rect 4905 16541 4939 16575
rect 9505 16541 9539 16575
rect 10701 16541 10735 16575
rect 12173 16541 12207 16575
rect 16129 16541 16163 16575
rect 16681 16541 16715 16575
rect 17785 16541 17819 16575
rect 23673 16541 23707 16575
rect 25145 16541 25179 16575
rect 28825 16541 28859 16575
rect 29745 16541 29779 16575
rect 2513 16473 2547 16507
rect 6009 16473 6043 16507
rect 8217 16473 8251 16507
rect 14381 16473 14415 16507
rect 15393 16473 15427 16507
rect 19717 16473 19751 16507
rect 21465 16473 21499 16507
rect 23029 16473 23063 16507
rect 27629 16473 27663 16507
rect 6653 16405 6687 16439
rect 7021 16405 7055 16439
rect 7849 16405 7883 16439
rect 9137 16405 9171 16439
rect 11345 16405 11379 16439
rect 13369 16405 13403 16439
rect 15025 16405 15059 16439
rect 15485 16405 15519 16439
rect 17325 16405 17359 16439
rect 18429 16405 18463 16439
rect 21925 16405 21959 16439
rect 22293 16405 22327 16439
rect 23765 16405 23799 16439
rect 24777 16405 24811 16439
rect 27261 16405 27295 16439
rect 28457 16405 28491 16439
rect 5641 16201 5675 16235
rect 5733 16201 5767 16235
rect 7849 16201 7883 16235
rect 8953 16201 8987 16235
rect 14841 16201 14875 16235
rect 16681 16201 16715 16235
rect 16957 16201 16991 16235
rect 17877 16201 17911 16235
rect 20085 16201 20119 16235
rect 22477 16201 22511 16235
rect 24133 16201 24167 16235
rect 4445 16133 4479 16167
rect 7113 16133 7147 16167
rect 9689 16133 9723 16167
rect 10517 16133 10551 16167
rect 11345 16133 11379 16167
rect 14013 16133 14047 16167
rect 18521 16133 18555 16167
rect 18705 16133 18739 16167
rect 24041 16133 24075 16167
rect 1777 16065 1811 16099
rect 3617 16065 3651 16099
rect 7021 16065 7055 16099
rect 8861 16065 8895 16099
rect 9873 16065 9907 16099
rect 11713 16065 11747 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 17049 16065 17083 16099
rect 17785 16065 17819 16099
rect 18981 16065 19015 16099
rect 20453 16065 20487 16099
rect 21465 16065 21499 16099
rect 22569 16065 22603 16099
rect 27169 16065 27203 16099
rect 28273 16065 28307 16099
rect 2053 15997 2087 16031
rect 5917 15997 5951 16031
rect 7297 15997 7331 16031
rect 9137 15997 9171 16031
rect 10609 15997 10643 16031
rect 10701 15997 10735 16031
rect 11989 15997 12023 16031
rect 14105 15997 14139 16031
rect 15117 15997 15151 16031
rect 18061 15997 18095 16031
rect 20545 15997 20579 16031
rect 20637 15997 20671 16031
rect 22661 15997 22695 16031
rect 23305 15997 23339 16031
rect 24317 15997 24351 16031
rect 24869 15997 24903 16031
rect 25145 15997 25179 16031
rect 27813 15997 27847 16031
rect 8493 15929 8527 15963
rect 10149 15929 10183 15963
rect 22109 15929 22143 15963
rect 23673 15929 23707 15963
rect 28917 15929 28951 15963
rect 5273 15861 5307 15895
rect 6653 15861 6687 15895
rect 13461 15861 13495 15895
rect 13829 15861 13863 15895
rect 14473 15861 14507 15895
rect 16313 15861 16347 15895
rect 17417 15861 17451 15895
rect 19625 15861 19659 15895
rect 21281 15861 21315 15895
rect 23213 15861 23247 15895
rect 26617 15861 26651 15895
rect 29561 15861 29595 15895
rect 7849 15657 7883 15691
rect 13277 15657 13311 15691
rect 14749 15657 14783 15691
rect 15945 15657 15979 15691
rect 18889 15657 18923 15691
rect 28641 15657 28675 15691
rect 5181 15589 5215 15623
rect 7481 15589 7515 15623
rect 20729 15589 20763 15623
rect 2053 15521 2087 15555
rect 4629 15521 4663 15555
rect 5825 15521 5859 15555
rect 6837 15521 6871 15555
rect 6929 15521 6963 15555
rect 8493 15521 8527 15555
rect 10149 15521 10183 15555
rect 10333 15521 10367 15555
rect 11529 15521 11563 15555
rect 12817 15521 12851 15555
rect 14473 15521 14507 15555
rect 15209 15521 15243 15555
rect 15393 15521 15427 15555
rect 16589 15521 16623 15555
rect 17141 15521 17175 15555
rect 19349 15521 19383 15555
rect 20177 15521 20211 15555
rect 20361 15521 20395 15555
rect 21097 15521 21131 15555
rect 23857 15521 23891 15555
rect 24593 15521 24627 15555
rect 25789 15521 25823 15555
rect 26893 15521 26927 15555
rect 26985 15521 27019 15555
rect 1777 15453 1811 15487
rect 4445 15453 4479 15487
rect 5549 15453 5583 15487
rect 6745 15453 6779 15487
rect 9229 15453 9263 15487
rect 10057 15453 10091 15487
rect 11345 15453 11379 15487
rect 12541 15453 12575 15487
rect 13737 15453 13771 15487
rect 16405 15453 16439 15487
rect 27629 15453 27663 15487
rect 5641 15385 5675 15419
rect 8309 15385 8343 15419
rect 9321 15385 9355 15419
rect 11437 15385 11471 15419
rect 15117 15385 15151 15419
rect 17417 15385 17451 15419
rect 21373 15385 21407 15419
rect 23673 15385 23707 15419
rect 25697 15385 25731 15419
rect 26801 15385 26835 15419
rect 3341 15317 3375 15351
rect 3525 15317 3559 15351
rect 3985 15317 4019 15351
rect 4353 15317 4387 15351
rect 6377 15317 6411 15351
rect 8217 15317 8251 15351
rect 8953 15317 8987 15351
rect 9689 15317 9723 15351
rect 10977 15317 11011 15351
rect 11989 15317 12023 15351
rect 12173 15317 12207 15351
rect 12633 15317 12667 15351
rect 13553 15317 13587 15351
rect 14197 15317 14231 15351
rect 16313 15317 16347 15351
rect 19717 15317 19751 15351
rect 20085 15317 20119 15351
rect 22845 15317 22879 15351
rect 23305 15317 23339 15351
rect 23765 15317 23799 15351
rect 25237 15317 25271 15351
rect 25605 15317 25639 15351
rect 26433 15317 26467 15351
rect 28273 15317 28307 15351
rect 4169 15113 4203 15147
rect 4997 15113 5031 15147
rect 12449 15113 12483 15147
rect 16313 15113 16347 15147
rect 17049 15113 17083 15147
rect 27445 15113 27479 15147
rect 27629 15113 27663 15147
rect 9965 15045 9999 15079
rect 14841 15045 14875 15079
rect 19993 15045 20027 15079
rect 23857 15045 23891 15079
rect 27721 15045 27755 15079
rect 1777 14977 1811 15011
rect 3525 14977 3559 15011
rect 6009 14977 6043 15011
rect 6837 14977 6871 15011
rect 7941 14977 7975 15011
rect 10793 14977 10827 15011
rect 11805 14977 11839 15011
rect 12817 14977 12851 15011
rect 12909 14977 12943 15011
rect 14105 14977 14139 15011
rect 14565 14977 14599 15011
rect 16865 14977 16899 15011
rect 17325 14977 17359 15011
rect 19717 14977 19751 15011
rect 22017 14977 22051 15011
rect 23121 14977 23155 15011
rect 27905 14977 27939 15011
rect 2053 14909 2087 14943
rect 5089 14909 5123 14943
rect 5273 14909 5307 14943
rect 8217 14909 8251 14943
rect 10885 14909 10919 14943
rect 10977 14909 11011 14943
rect 13001 14909 13035 14943
rect 21465 14909 21499 14943
rect 24869 14909 24903 14943
rect 25145 14909 25179 14943
rect 6561 14841 6595 14875
rect 13921 14841 13955 14875
rect 18613 14841 18647 14875
rect 27261 14841 27295 14875
rect 4629 14773 4663 14807
rect 5825 14773 5859 14807
rect 7481 14773 7515 14807
rect 10425 14773 10459 14807
rect 11897 14773 11931 14807
rect 13553 14773 13587 14807
rect 19441 14773 19475 14807
rect 22661 14773 22695 14807
rect 24317 14773 24351 14807
rect 24593 14773 24627 14807
rect 26617 14773 26651 14807
rect 27077 14773 27111 14807
rect 4169 14569 4203 14603
rect 9413 14569 9447 14603
rect 11713 14569 11747 14603
rect 13737 14569 13771 14603
rect 14197 14569 14231 14603
rect 18613 14569 18647 14603
rect 18981 14569 19015 14603
rect 21925 14569 21959 14603
rect 24041 14569 24075 14603
rect 27169 14569 27203 14603
rect 2053 14433 2087 14467
rect 3617 14433 3651 14467
rect 4813 14433 4847 14467
rect 5641 14433 5675 14467
rect 7389 14433 7423 14467
rect 8309 14433 8343 14467
rect 8401 14433 8435 14467
rect 9873 14433 9907 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 14933 14433 14967 14467
rect 17141 14433 17175 14467
rect 19993 14433 20027 14467
rect 21189 14433 21223 14467
rect 22293 14433 22327 14467
rect 1777 14365 1811 14399
rect 5365 14365 5399 14399
rect 9781 14365 9815 14399
rect 11069 14365 11103 14399
rect 11989 14365 12023 14399
rect 14657 14365 14691 14399
rect 16865 14365 16899 14399
rect 19901 14365 19935 14399
rect 26525 14365 26559 14399
rect 12265 14297 12299 14331
rect 21005 14297 21039 14331
rect 21741 14297 21775 14331
rect 22569 14297 22603 14331
rect 24869 14297 24903 14331
rect 25145 14297 25179 14331
rect 25973 14297 26007 14331
rect 3341 14229 3375 14263
rect 3801 14229 3835 14263
rect 4537 14229 4571 14263
rect 4629 14229 4663 14263
rect 7849 14229 7883 14263
rect 8217 14229 8251 14263
rect 9045 14229 9079 14263
rect 10609 14229 10643 14263
rect 10977 14229 11011 14263
rect 16405 14229 16439 14263
rect 19441 14229 19475 14263
rect 19809 14229 19843 14263
rect 20637 14229 20671 14263
rect 21097 14229 21131 14263
rect 24409 14229 24443 14263
rect 24685 14229 24719 14263
rect 3525 14025 3559 14059
rect 6469 14025 6503 14059
rect 7297 14025 7331 14059
rect 8125 14025 8159 14059
rect 8493 14025 8527 14059
rect 8585 14025 8619 14059
rect 11069 14025 11103 14059
rect 13093 14025 13127 14059
rect 13369 14025 13403 14059
rect 14565 14025 14599 14059
rect 15393 14025 15427 14059
rect 15853 14025 15887 14059
rect 16405 14025 16439 14059
rect 18889 14025 18923 14059
rect 19257 14025 19291 14059
rect 19533 14025 19567 14059
rect 21373 14025 21407 14059
rect 21557 14025 21591 14059
rect 22477 14025 22511 14059
rect 23213 14025 23247 14059
rect 24409 14025 24443 14059
rect 25513 14025 25547 14059
rect 26249 14025 26283 14059
rect 26709 14025 26743 14059
rect 7389 13957 7423 13991
rect 15761 13957 15795 13991
rect 16773 13957 16807 13991
rect 23673 13957 23707 13991
rect 25421 13957 25455 13991
rect 26065 13957 26099 13991
rect 1777 13889 1811 13923
rect 3709 13889 3743 13923
rect 4169 13889 4203 13923
rect 11713 13889 11747 13923
rect 11989 13889 12023 13923
rect 14473 13889 14507 13923
rect 17141 13889 17175 13923
rect 20545 13889 20579 13923
rect 20637 13889 20671 13923
rect 22385 13889 22419 13923
rect 23581 13889 23615 13923
rect 24593 13889 24627 13923
rect 26525 13889 26559 13923
rect 2053 13821 2087 13855
rect 4445 13821 4479 13855
rect 5917 13821 5951 13855
rect 6653 13821 6687 13855
rect 7573 13821 7607 13855
rect 8769 13821 8803 13855
rect 9321 13821 9355 13855
rect 9597 13821 9631 13855
rect 12909 13821 12943 13855
rect 13277 13821 13311 13855
rect 13553 13821 13587 13855
rect 14749 13821 14783 13855
rect 15945 13821 15979 13855
rect 17417 13821 17451 13855
rect 20821 13821 20855 13855
rect 21189 13821 21223 13855
rect 22569 13821 22603 13855
rect 23765 13821 23799 13855
rect 25697 13821 25731 13855
rect 13829 13753 13863 13787
rect 14105 13753 14139 13787
rect 20177 13753 20211 13787
rect 6929 13685 6963 13719
rect 22017 13685 22051 13719
rect 25053 13685 25087 13719
rect 3617 13481 3651 13515
rect 14546 13481 14580 13515
rect 16037 13481 16071 13515
rect 22017 13481 22051 13515
rect 22937 13481 22971 13515
rect 3433 13413 3467 13447
rect 4445 13413 4479 13447
rect 8585 13413 8619 13447
rect 11437 13413 11471 13447
rect 11621 13413 11655 13447
rect 13737 13413 13771 13447
rect 18889 13413 18923 13447
rect 24593 13413 24627 13447
rect 2053 13345 2087 13379
rect 4905 13345 4939 13379
rect 4997 13345 5031 13379
rect 6193 13345 6227 13379
rect 7113 13345 7147 13379
rect 9781 13345 9815 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 17141 13345 17175 13379
rect 20545 13345 20579 13379
rect 23765 13345 23799 13379
rect 23857 13345 23891 13379
rect 25145 13345 25179 13379
rect 1777 13277 1811 13311
rect 4813 13277 4847 13311
rect 6101 13277 6135 13311
rect 6837 13277 6871 13311
rect 10793 13277 10827 13311
rect 19901 13277 19935 13311
rect 20269 13277 20303 13311
rect 22661 13277 22695 13311
rect 23673 13277 23707 13311
rect 24961 13277 24995 13311
rect 25789 13277 25823 13311
rect 3985 13209 4019 13243
rect 10701 13209 10735 13243
rect 12265 13209 12299 13243
rect 17417 13209 17451 13243
rect 4169 13141 4203 13175
rect 5641 13141 5675 13175
rect 6009 13141 6043 13175
rect 9137 13141 9171 13175
rect 9505 13141 9539 13175
rect 9597 13141 9631 13175
rect 10333 13141 10367 13175
rect 19441 13141 19475 13175
rect 22477 13141 22511 13175
rect 23305 13141 23339 13175
rect 25053 13141 25087 13175
rect 26433 13141 26467 13175
rect 2881 12937 2915 12971
rect 7297 12937 7331 12971
rect 11897 12937 11931 12971
rect 12817 12937 12851 12971
rect 14381 12937 14415 12971
rect 15577 12937 15611 12971
rect 16037 12937 16071 12971
rect 17141 12937 17175 12971
rect 17509 12937 17543 12971
rect 17601 12937 17635 12971
rect 18705 12937 18739 12971
rect 3801 12869 3835 12903
rect 6377 12869 6411 12903
rect 10149 12869 10183 12903
rect 10517 12869 10551 12903
rect 14749 12869 14783 12903
rect 19533 12869 19567 12903
rect 20269 12869 20303 12903
rect 20913 12869 20947 12903
rect 21649 12869 21683 12903
rect 1593 12801 1627 12835
rect 3157 12801 3191 12835
rect 4261 12801 4295 12835
rect 7389 12801 7423 12835
rect 8125 12801 8159 12835
rect 10609 12801 10643 12835
rect 10793 12801 10827 12835
rect 13461 12801 13495 12835
rect 14105 12801 14139 12835
rect 15945 12801 15979 12835
rect 22477 12801 22511 12835
rect 25237 12801 25271 12835
rect 1869 12733 1903 12767
rect 4537 12733 4571 12767
rect 6009 12733 6043 12767
rect 7573 12733 7607 12767
rect 8401 12733 8435 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 12909 12733 12943 12767
rect 13093 12733 13127 12767
rect 14841 12733 14875 12767
rect 15025 12733 15059 12767
rect 16221 12733 16255 12767
rect 16681 12733 16715 12767
rect 17693 12733 17727 12767
rect 18797 12733 18831 12767
rect 18981 12733 19015 12767
rect 22017 12733 22051 12767
rect 23029 12733 23063 12767
rect 23305 12733 23339 12767
rect 6929 12665 6963 12699
rect 11529 12665 11563 12699
rect 6561 12597 6595 12631
rect 12081 12597 12115 12631
rect 12449 12597 12483 12631
rect 13737 12597 13771 12631
rect 13829 12597 13863 12631
rect 18337 12597 18371 12631
rect 24777 12597 24811 12631
rect 25881 12597 25915 12631
rect 2329 12393 2363 12427
rect 4169 12393 4203 12427
rect 5089 12393 5123 12427
rect 14473 12393 14507 12427
rect 17969 12393 18003 12427
rect 14105 12325 14139 12359
rect 18613 12325 18647 12359
rect 24593 12325 24627 12359
rect 5549 12257 5583 12291
rect 5825 12257 5859 12291
rect 7573 12257 7607 12291
rect 8401 12257 8435 12291
rect 9873 12257 9907 12291
rect 11161 12257 11195 12291
rect 12449 12257 12483 12291
rect 13645 12257 13679 12291
rect 15577 12257 15611 12291
rect 16221 12257 16255 12291
rect 20361 12257 20395 12291
rect 22293 12257 22327 12291
rect 25053 12257 25087 12291
rect 25145 12257 25179 12291
rect 1685 12189 1719 12223
rect 2789 12189 2823 12223
rect 3433 12189 3467 12223
rect 4445 12189 4479 12223
rect 9137 12189 9171 12223
rect 12173 12189 12207 12223
rect 13461 12189 13495 12223
rect 14841 12189 14875 12223
rect 18797 12189 18831 12223
rect 19625 12189 19659 12223
rect 20085 12189 20119 12223
rect 24961 12189 24995 12223
rect 11069 12121 11103 12155
rect 12265 12121 12299 12155
rect 16497 12121 16531 12155
rect 22569 12121 22603 12155
rect 3985 12053 4019 12087
rect 7849 12053 7883 12087
rect 8033 12053 8067 12087
rect 10609 12053 10643 12087
rect 10977 12053 11011 12087
rect 11805 12053 11839 12087
rect 13001 12053 13035 12087
rect 13369 12053 13403 12087
rect 14381 12053 14415 12087
rect 18245 12053 18279 12087
rect 19349 12053 19383 12087
rect 19441 12053 19475 12087
rect 21833 12053 21867 12087
rect 24041 12053 24075 12087
rect 25605 12053 25639 12087
rect 2329 11849 2363 11883
rect 2789 11849 2823 11883
rect 3709 11849 3743 11883
rect 4813 11849 4847 11883
rect 5641 11849 5675 11883
rect 6745 11849 6779 11883
rect 10977 11849 11011 11883
rect 12449 11849 12483 11883
rect 16773 11849 16807 11883
rect 17693 11849 17727 11883
rect 9597 11781 9631 11815
rect 12357 11781 12391 11815
rect 13461 11781 13495 11815
rect 21925 11781 21959 11815
rect 1685 11713 1719 11747
rect 3065 11713 3099 11747
rect 4169 11713 4203 11747
rect 5733 11713 5767 11747
rect 6653 11713 6687 11747
rect 11621 11713 11655 11747
rect 13185 11713 13219 11747
rect 15393 11713 15427 11747
rect 17601 11713 17635 11747
rect 18429 11713 18463 11747
rect 18705 11713 18739 11747
rect 22385 11713 22419 11747
rect 5825 11645 5859 11679
rect 7389 11645 7423 11679
rect 7665 11645 7699 11679
rect 10333 11645 10367 11679
rect 12633 11645 12667 11679
rect 16221 11645 16255 11679
rect 16957 11645 16991 11679
rect 17785 11645 17819 11679
rect 19717 11645 19751 11679
rect 19993 11645 20027 11679
rect 22661 11645 22695 11679
rect 11989 11577 12023 11611
rect 17233 11577 17267 11611
rect 5273 11509 5307 11543
rect 9137 11509 9171 11543
rect 14933 11509 14967 11543
rect 21465 11509 21499 11543
rect 24133 11509 24167 11543
rect 24409 11509 24443 11543
rect 24593 11509 24627 11543
rect 2881 11305 2915 11339
rect 4169 11305 4203 11339
rect 7205 11305 7239 11339
rect 7849 11305 7883 11339
rect 9229 11305 9263 11339
rect 10425 11305 10459 11339
rect 13737 11305 13771 11339
rect 14197 11305 14231 11339
rect 16589 11305 16623 11339
rect 23765 11305 23799 11339
rect 3433 11237 3467 11271
rect 18889 11237 18923 11271
rect 22661 11237 22695 11271
rect 1869 11169 1903 11203
rect 4997 11169 5031 11203
rect 8401 11169 8435 11203
rect 9781 11169 9815 11203
rect 11069 11169 11103 11203
rect 13369 11169 13403 11203
rect 14841 11169 14875 11203
rect 17417 11169 17451 11203
rect 29745 11169 29779 11203
rect 1501 11101 1535 11135
rect 1593 11101 1627 11135
rect 3249 11101 3283 11135
rect 4077 11101 4111 11135
rect 7389 11101 7423 11135
rect 8309 11101 8343 11135
rect 9597 11101 9631 11135
rect 10793 11101 10827 11135
rect 11621 11101 11655 11135
rect 13921 11101 13955 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 17141 11101 17175 11135
rect 20361 11101 20395 11135
rect 20913 11101 20947 11135
rect 23121 11101 23155 11135
rect 32045 11101 32079 11135
rect 5273 11033 5307 11067
rect 10333 11033 10367 11067
rect 10885 11033 10919 11067
rect 11897 11033 11931 11067
rect 15117 11033 15151 11067
rect 19533 11033 19567 11067
rect 21189 11033 21223 11067
rect 24133 11033 24167 11067
rect 30021 11033 30055 11067
rect 31769 11033 31803 11067
rect 4629 10965 4663 10999
rect 6745 10965 6779 10999
rect 8217 10965 8251 10999
rect 9689 10965 9723 10999
rect 1501 10761 1535 10795
rect 1777 10761 1811 10795
rect 3433 10761 3467 10795
rect 3801 10761 3835 10795
rect 4905 10761 4939 10795
rect 6009 10761 6043 10795
rect 6929 10761 6963 10795
rect 10149 10761 10183 10795
rect 11621 10761 11655 10795
rect 11805 10761 11839 10795
rect 14381 10761 14415 10795
rect 14841 10761 14875 10795
rect 16865 10761 16899 10795
rect 21465 10761 21499 10795
rect 21833 10761 21867 10795
rect 22845 10761 22879 10795
rect 2329 10693 2363 10727
rect 3893 10693 3927 10727
rect 10793 10693 10827 10727
rect 15945 10693 15979 10727
rect 16037 10693 16071 10727
rect 2145 10625 2179 10659
rect 2789 10625 2823 10659
rect 4261 10625 4295 10659
rect 5365 10625 5399 10659
rect 12173 10625 12207 10659
rect 14749 10625 14783 10659
rect 17509 10625 17543 10659
rect 22201 10625 22235 10659
rect 23305 10625 23339 10659
rect 7021 10557 7055 10591
rect 7113 10557 7147 10591
rect 7757 10557 7791 10591
rect 8033 10557 8067 10591
rect 9781 10557 9815 10591
rect 10885 10557 10919 10591
rect 10977 10557 11011 10591
rect 12449 10557 12483 10591
rect 15025 10557 15059 10591
rect 16221 10557 16255 10591
rect 17785 10557 17819 10591
rect 19717 10557 19751 10591
rect 19993 10557 20027 10591
rect 23949 10557 23983 10591
rect 15577 10489 15611 10523
rect 6561 10421 6595 10455
rect 10425 10421 10459 10455
rect 13921 10421 13955 10455
rect 19257 10421 19291 10455
rect 3065 10217 3099 10251
rect 3617 10217 3651 10251
rect 4169 10217 4203 10251
rect 6193 10217 6227 10251
rect 6653 10217 6687 10251
rect 13645 10217 13679 10251
rect 16681 10217 16715 10251
rect 18889 10217 18923 10251
rect 22385 10217 22419 10251
rect 13921 10149 13955 10183
rect 16405 10149 16439 10183
rect 1593 10081 1627 10115
rect 7205 10081 7239 10115
rect 8309 10081 8343 10115
rect 8401 10081 8435 10115
rect 14657 10081 14691 10115
rect 17141 10081 17175 10115
rect 19533 10081 19567 10115
rect 19809 10081 19843 10115
rect 1869 10013 1903 10047
rect 4997 10013 5031 10047
rect 5549 10013 5583 10047
rect 7113 10013 7147 10047
rect 9137 10013 9171 10047
rect 11437 10013 11471 10047
rect 21741 10013 21775 10047
rect 2973 9945 3007 9979
rect 4077 9945 4111 9979
rect 4813 9945 4847 9979
rect 9413 9945 9447 9979
rect 11713 9945 11747 9979
rect 14933 9945 14967 9979
rect 17417 9945 17451 9979
rect 7021 9877 7055 9911
rect 7849 9877 7883 9911
rect 8217 9877 8251 9911
rect 10885 9877 10919 9911
rect 13185 9877 13219 9911
rect 13461 9877 13495 9911
rect 14105 9877 14139 9911
rect 14289 9877 14323 9911
rect 21281 9877 21315 9911
rect 21373 9673 21407 9707
rect 21557 9673 21591 9707
rect 1501 9605 1535 9639
rect 1777 9605 1811 9639
rect 3341 9605 3375 9639
rect 6009 9605 6043 9639
rect 7941 9605 7975 9639
rect 8677 9605 8711 9639
rect 10701 9605 10735 9639
rect 13737 9605 13771 9639
rect 17141 9605 17175 9639
rect 19533 9605 19567 9639
rect 20913 9605 20947 9639
rect 22661 9605 22695 9639
rect 27813 9605 27847 9639
rect 2421 9537 2455 9571
rect 4077 9537 4111 9571
rect 5365 9537 5399 9571
rect 7297 9537 7331 9571
rect 10425 9537 10459 9571
rect 10977 9537 11011 9571
rect 11713 9537 11747 9571
rect 14565 9537 14599 9571
rect 16865 9537 16899 9571
rect 19441 9537 19475 9571
rect 20269 9537 20303 9571
rect 22017 9537 22051 9571
rect 27169 9537 27203 9571
rect 2145 9469 2179 9503
rect 3709 9469 3743 9503
rect 4261 9469 4295 9503
rect 4721 9469 4755 9503
rect 6653 9469 6687 9503
rect 8401 9469 8435 9503
rect 11989 9469 12023 9503
rect 13461 9469 13495 9503
rect 14013 9469 14047 9503
rect 14841 9469 14875 9503
rect 16313 9469 16347 9503
rect 19717 9469 19751 9503
rect 3433 9401 3467 9435
rect 19073 9401 19107 9435
rect 1685 9333 1719 9367
rect 3893 9333 3927 9367
rect 4629 9333 4663 9367
rect 10149 9333 10183 9367
rect 14197 9333 14231 9367
rect 18613 9333 18647 9367
rect 1593 9129 1627 9163
rect 2053 9129 2087 9163
rect 4721 9129 4755 9163
rect 4997 9129 5031 9163
rect 6285 9129 6319 9163
rect 7389 9129 7423 9163
rect 10425 9129 10459 9163
rect 18889 9129 18923 9163
rect 19441 9129 19475 9163
rect 21005 9129 21039 9163
rect 27905 9129 27939 9163
rect 28733 9129 28767 9163
rect 9965 9061 9999 9095
rect 14381 9061 14415 9095
rect 15669 9061 15703 9095
rect 2605 8993 2639 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 10977 8993 11011 9027
rect 12173 8993 12207 9027
rect 12909 8993 12943 9027
rect 13185 8993 13219 9027
rect 15025 8993 15059 9027
rect 16037 8993 16071 9027
rect 1777 8925 1811 8959
rect 2881 8925 2915 8959
rect 4077 8925 4111 8959
rect 5181 8925 5215 8959
rect 5641 8925 5675 8959
rect 6745 8925 6779 8959
rect 8217 8925 8251 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 10885 8925 10919 8959
rect 18245 8925 18279 8959
rect 20361 8925 20395 8959
rect 27629 8925 27663 8959
rect 4261 8857 4295 8891
rect 11989 8857 12023 8891
rect 12081 8857 12115 8891
rect 14841 8857 14875 8891
rect 16313 8857 16347 8891
rect 2329 8789 2363 8823
rect 7849 8789 7883 8823
rect 10793 8789 10827 8823
rect 11621 8789 11655 8823
rect 14749 8789 14783 8823
rect 17785 8789 17819 8823
rect 19533 8789 19567 8823
rect 19717 8789 19751 8823
rect 19901 8789 19935 8823
rect 28089 8789 28123 8823
rect 28549 8789 28583 8823
rect 1593 8585 1627 8619
rect 5181 8585 5215 8619
rect 5733 8585 5767 8619
rect 5825 8585 5859 8619
rect 9873 8585 9907 8619
rect 10241 8585 10275 8619
rect 11069 8585 11103 8619
rect 11345 8585 11379 8619
rect 11621 8585 11655 8619
rect 11897 8585 11931 8619
rect 14381 8585 14415 8619
rect 16313 8585 16347 8619
rect 17877 8585 17911 8619
rect 18245 8585 18279 8619
rect 19257 8585 19291 8619
rect 9413 8517 9447 8551
rect 10333 8517 10367 8551
rect 12265 8517 12299 8551
rect 14841 8517 14875 8551
rect 1777 8449 1811 8483
rect 2329 8449 2363 8483
rect 3617 8449 3651 8483
rect 6561 8449 6595 8483
rect 7941 8449 7975 8483
rect 8493 8449 8527 8483
rect 8769 8449 8803 8483
rect 12357 8449 12391 8483
rect 13461 8449 13495 8483
rect 14749 8449 14783 8483
rect 15669 8449 15703 8483
rect 17233 8449 17267 8483
rect 18613 8449 18647 8483
rect 2053 8381 2087 8415
rect 3341 8381 3375 8415
rect 4537 8381 4571 8415
rect 4629 8381 4663 8415
rect 6837 8381 6871 8415
rect 8125 8381 8159 8415
rect 10517 8381 10551 8415
rect 12541 8381 12575 8415
rect 13553 8381 13587 8415
rect 13737 8381 13771 8415
rect 14933 8381 14967 8415
rect 16681 8381 16715 8415
rect 10977 8313 11011 8347
rect 13093 8313 13127 8347
rect 19533 8313 19567 8347
rect 5365 8245 5399 8279
rect 5457 8245 5491 8279
rect 1593 8041 1627 8075
rect 5365 8041 5399 8075
rect 8585 8041 8619 8075
rect 11161 8041 11195 8075
rect 12357 8041 12391 8075
rect 13461 8041 13495 8075
rect 14289 8041 14323 8075
rect 16773 8041 16807 8075
rect 18797 8041 18831 8075
rect 3985 7973 4019 8007
rect 10149 7973 10183 8007
rect 17233 7973 17267 8007
rect 2237 7905 2271 7939
rect 2881 7905 2915 7939
rect 7205 7905 7239 7939
rect 9413 7905 9447 7939
rect 10609 7905 10643 7939
rect 10793 7905 10827 7939
rect 14749 7905 14783 7939
rect 14933 7905 14967 7939
rect 1777 7837 1811 7871
rect 4169 7837 4203 7871
rect 4905 7837 4939 7871
rect 5273 7837 5307 7871
rect 5917 7837 5951 7871
rect 6193 7837 6227 7871
rect 7941 7837 7975 7871
rect 9229 7837 9263 7871
rect 10517 7837 10551 7871
rect 11713 7837 11747 7871
rect 12817 7837 12851 7871
rect 15485 7837 15519 7871
rect 16129 7837 16163 7871
rect 17417 7837 17451 7871
rect 18153 7837 18187 7871
rect 3525 7769 3559 7803
rect 3341 7701 3375 7735
rect 4721 7701 4755 7735
rect 5641 7701 5675 7735
rect 9873 7701 9907 7735
rect 11345 7701 11379 7735
rect 14657 7701 14691 7735
rect 2789 7497 2823 7531
rect 4537 7497 4571 7531
rect 4721 7497 4755 7531
rect 4905 7497 4939 7531
rect 5825 7497 5859 7531
rect 7113 7497 7147 7531
rect 7941 7497 7975 7531
rect 9597 7497 9631 7531
rect 11253 7497 11287 7531
rect 11805 7497 11839 7531
rect 13737 7497 13771 7531
rect 16037 7497 16071 7531
rect 24041 7497 24075 7531
rect 16865 7429 16899 7463
rect 1869 7361 1903 7395
rect 3617 7361 3651 7395
rect 6009 7361 6043 7395
rect 6653 7361 6687 7395
rect 7389 7361 7423 7395
rect 8309 7361 8343 7395
rect 10609 7361 10643 7395
rect 11989 7361 12023 7395
rect 13093 7361 13127 7395
rect 14289 7361 14323 7395
rect 15393 7361 15427 7395
rect 22293 7361 22327 7395
rect 24317 7361 24351 7395
rect 1593 7293 1627 7327
rect 2881 7293 2915 7327
rect 3341 7293 3375 7327
rect 5181 7293 5215 7327
rect 6837 7293 6871 7327
rect 8585 7293 8619 7327
rect 10701 7293 10735 7327
rect 10885 7293 10919 7327
rect 14933 7293 14967 7327
rect 22569 7293 22603 7327
rect 7481 7225 7515 7259
rect 10241 7225 10275 7259
rect 7757 7157 7791 7191
rect 12357 7157 12391 7191
rect 12541 7157 12575 7191
rect 7205 6953 7239 6987
rect 1869 6817 1903 6851
rect 2697 6817 2731 6851
rect 2881 6817 2915 6851
rect 3985 6817 4019 6851
rect 7665 6817 7699 6851
rect 10333 6817 10367 6851
rect 12173 6817 12207 6851
rect 21373 6817 21407 6851
rect 1593 6749 1627 6783
rect 4905 6749 4939 6783
rect 5365 6749 5399 6783
rect 6009 6749 6043 6783
rect 6653 6749 6687 6783
rect 7941 6749 7975 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 11529 6749 11563 6783
rect 12633 6749 12667 6783
rect 14289 6749 14323 6783
rect 15117 6749 15151 6783
rect 20729 6749 20763 6783
rect 3341 6681 3375 6715
rect 4169 6681 4203 6715
rect 4261 6681 4295 6715
rect 7389 6681 7423 6715
rect 10517 6681 10551 6715
rect 10885 6681 10919 6715
rect 11069 6681 11103 6715
rect 13277 6681 13311 6715
rect 5181 6613 5215 6647
rect 5825 6613 5859 6647
rect 6469 6613 6503 6647
rect 7021 6613 7055 6647
rect 14933 6613 14967 6647
rect 2789 6409 2823 6443
rect 3065 6409 3099 6443
rect 3985 6409 4019 6443
rect 4629 6409 4663 6443
rect 5825 6409 5859 6443
rect 6193 6409 6227 6443
rect 8677 6409 8711 6443
rect 9597 6409 9631 6443
rect 12173 6409 12207 6443
rect 14289 6409 14323 6443
rect 23949 6341 23983 6375
rect 1593 6273 1627 6307
rect 1869 6273 1903 6307
rect 3525 6273 3559 6307
rect 4169 6273 4203 6307
rect 5457 6273 5491 6307
rect 5917 6273 5951 6307
rect 10333 6273 10367 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 12909 6273 12943 6307
rect 23029 6273 23063 6307
rect 6929 6205 6963 6239
rect 8861 6205 8895 6239
rect 8953 6205 8987 6239
rect 13553 6205 13587 6239
rect 3341 6137 3375 6171
rect 5273 6069 5307 6103
rect 23305 6069 23339 6103
rect 23489 6069 23523 6103
rect 2881 5865 2915 5899
rect 3985 5865 4019 5899
rect 5273 5865 5307 5899
rect 9137 5865 9171 5899
rect 9689 5865 9723 5899
rect 11713 5865 11747 5899
rect 19349 5865 19383 5899
rect 22845 5865 22879 5899
rect 1869 5729 1903 5763
rect 3341 5729 3375 5763
rect 5733 5729 5767 5763
rect 14841 5729 14875 5763
rect 17141 5729 17175 5763
rect 18889 5729 18923 5763
rect 25973 5729 26007 5763
rect 26709 5729 26743 5763
rect 1593 5661 1627 5695
rect 3065 5661 3099 5695
rect 3617 5661 3651 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 5457 5661 5491 5695
rect 9321 5661 9355 5695
rect 11897 5661 11931 5695
rect 13645 5661 13679 5695
rect 14381 5661 14415 5695
rect 22344 5661 22378 5695
rect 25789 5661 25823 5695
rect 14565 5593 14599 5627
rect 17417 5593 17451 5627
rect 22431 5593 22465 5627
rect 4629 5525 4663 5559
rect 12817 5525 12851 5559
rect 13461 5525 13495 5559
rect 16589 5525 16623 5559
rect 4169 5321 4203 5355
rect 22431 5321 22465 5355
rect 4905 5253 4939 5287
rect 24961 5253 24995 5287
rect 26617 5253 26651 5287
rect 29009 5253 29043 5287
rect 1869 5185 1903 5219
rect 3065 5185 3099 5219
rect 3709 5185 3743 5219
rect 4353 5185 4387 5219
rect 4629 5185 4663 5219
rect 20913 5185 20947 5219
rect 21833 5185 21867 5219
rect 22360 5185 22394 5219
rect 1593 5117 1627 5151
rect 4997 5117 5031 5151
rect 24777 5117 24811 5151
rect 27169 5117 27203 5151
rect 27353 5117 27387 5151
rect 29469 5117 29503 5151
rect 29653 5117 29687 5151
rect 31309 5117 31343 5151
rect 3525 5049 3559 5083
rect 21373 5049 21407 5083
rect 2881 4981 2915 5015
rect 21005 4981 21039 5015
rect 2881 4777 2915 4811
rect 3433 4777 3467 4811
rect 3617 4777 3651 4811
rect 14933 4777 14967 4811
rect 19533 4777 19567 4811
rect 23075 4777 23109 4811
rect 3985 4709 4019 4743
rect 24731 4709 24765 4743
rect 1593 4641 1627 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 15761 4641 15795 4675
rect 17417 4641 17451 4675
rect 1869 4573 1903 4607
rect 3065 4573 3099 4607
rect 4169 4573 4203 4607
rect 4445 4573 4479 4607
rect 14289 4573 14323 4607
rect 19441 4573 19475 4607
rect 20269 4573 20303 4607
rect 22972 4573 23006 4607
rect 24628 4573 24662 4607
rect 15945 4505 15979 4539
rect 19901 4437 19935 4471
rect 1593 4097 1627 4131
rect 1869 4097 1903 4131
rect 3065 4097 3099 4131
rect 3709 4097 3743 4131
rect 3985 4097 4019 4131
rect 16865 4097 16899 4131
rect 4169 4029 4203 4063
rect 17049 4029 17083 4063
rect 18705 4029 18739 4063
rect 2881 3961 2915 3995
rect 3525 3961 3559 3995
rect 3525 3689 3559 3723
rect 3985 3689 4019 3723
rect 12173 3689 12207 3723
rect 2881 3621 2915 3655
rect 3433 3621 3467 3655
rect 1593 3553 1627 3587
rect 4629 3553 4663 3587
rect 1869 3485 1903 3519
rect 3065 3485 3099 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 2881 3145 2915 3179
rect 3525 3145 3559 3179
rect 10609 3145 10643 3179
rect 12725 3145 12759 3179
rect 11805 3077 11839 3111
rect 12633 3077 12667 3111
rect 14105 3077 14139 3111
rect 15853 3077 15887 3111
rect 18705 3077 18739 3111
rect 3065 3009 3099 3043
rect 3709 3009 3743 3043
rect 3985 3009 4019 3043
rect 8861 3009 8895 3043
rect 10885 3009 10919 3043
rect 18521 3009 18555 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 9137 2941 9171 2975
rect 14289 2941 14323 2975
rect 20361 2941 20395 2975
rect 4169 2873 4203 2907
rect 4353 2805 4387 2839
rect 11897 2805 11931 2839
rect 15945 2805 15979 2839
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 1593 2465 1627 2499
rect 1869 2465 1903 2499
rect 3525 2465 3559 2499
rect 4629 2465 4663 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 36369 2465 36403 2499
rect 3065 2397 3099 2431
rect 3801 2397 3835 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 25697 2397 25731 2431
rect 25973 2397 26007 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33701 2397 33735 2431
rect 33977 2397 34011 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 2881 2261 2915 2295
rect 3341 2261 3375 2295
<< metal1 >>
rect 8846 26120 8852 26172
rect 8904 26160 8910 26172
rect 30926 26160 30932 26172
rect 8904 26132 30932 26160
rect 8904 26120 8910 26132
rect 30926 26120 30932 26132
rect 30984 26120 30990 26172
rect 17862 26052 17868 26104
rect 17920 26092 17926 26104
rect 33962 26092 33968 26104
rect 17920 26064 33968 26092
rect 17920 26052 17926 26064
rect 33962 26052 33968 26064
rect 34020 26052 34026 26104
rect 15010 25984 15016 26036
rect 15068 26024 15074 26036
rect 35250 26024 35256 26036
rect 15068 25996 35256 26024
rect 15068 25984 15074 25996
rect 35250 25984 35256 25996
rect 35308 25984 35314 26036
rect 12434 25916 12440 25968
rect 12492 25956 12498 25968
rect 36078 25956 36084 25968
rect 12492 25928 36084 25956
rect 12492 25916 12498 25928
rect 36078 25916 36084 25928
rect 36136 25916 36142 25968
rect 17402 25848 17408 25900
rect 17460 25888 17466 25900
rect 40402 25888 40408 25900
rect 17460 25860 40408 25888
rect 17460 25848 17466 25860
rect 40402 25848 40408 25860
rect 40460 25848 40466 25900
rect 25038 25780 25044 25832
rect 25096 25820 25102 25832
rect 39758 25820 39764 25832
rect 25096 25792 39764 25820
rect 25096 25780 25102 25792
rect 39758 25780 39764 25792
rect 39816 25780 39822 25832
rect 11790 25712 11796 25764
rect 11848 25752 11854 25764
rect 36538 25752 36544 25764
rect 11848 25724 36544 25752
rect 11848 25712 11854 25724
rect 36538 25712 36544 25724
rect 36596 25712 36602 25764
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 38654 25684 38660 25696
rect 12308 25656 38660 25684
rect 12308 25644 12314 25656
rect 38654 25644 38660 25656
rect 38712 25644 38718 25696
rect 16666 25576 16672 25628
rect 16724 25616 16730 25628
rect 36262 25616 36268 25628
rect 16724 25588 36268 25616
rect 16724 25576 16730 25588
rect 36262 25576 36268 25588
rect 36320 25576 36326 25628
rect 6270 25508 6276 25560
rect 6328 25548 6334 25560
rect 35894 25548 35900 25560
rect 6328 25520 35900 25548
rect 6328 25508 6334 25520
rect 35894 25508 35900 25520
rect 35952 25508 35958 25560
rect 13538 25440 13544 25492
rect 13596 25480 13602 25492
rect 33318 25480 33324 25492
rect 13596 25452 33324 25480
rect 13596 25440 13602 25452
rect 33318 25440 33324 25452
rect 33376 25440 33382 25492
rect 11054 25372 11060 25424
rect 11112 25412 11118 25424
rect 34698 25412 34704 25424
rect 11112 25384 34704 25412
rect 11112 25372 11118 25384
rect 34698 25372 34704 25384
rect 34756 25372 34762 25424
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 34606 25344 34612 25356
rect 12124 25316 34612 25344
rect 12124 25304 12130 25316
rect 34606 25304 34612 25316
rect 34664 25304 34670 25356
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 32398 25276 32404 25288
rect 9916 25248 32404 25276
rect 9916 25236 9922 25248
rect 32398 25236 32404 25248
rect 32456 25236 32462 25288
rect 3878 25168 3884 25220
rect 3936 25208 3942 25220
rect 9766 25208 9772 25220
rect 3936 25180 9772 25208
rect 3936 25168 3942 25180
rect 9766 25168 9772 25180
rect 9824 25168 9830 25220
rect 22554 25168 22560 25220
rect 22612 25208 22618 25220
rect 32766 25208 32772 25220
rect 22612 25180 32772 25208
rect 22612 25168 22618 25180
rect 32766 25168 32772 25180
rect 32824 25168 32830 25220
rect 20622 25100 20628 25152
rect 20680 25140 20686 25152
rect 32674 25140 32680 25152
rect 20680 25112 32680 25140
rect 20680 25100 20686 25112
rect 32674 25100 32680 25112
rect 32732 25100 32738 25152
rect 6638 25032 6644 25084
rect 6696 25072 6702 25084
rect 22002 25072 22008 25084
rect 6696 25044 22008 25072
rect 6696 25032 6702 25044
rect 22002 25032 22008 25044
rect 22060 25032 22066 25084
rect 26142 25032 26148 25084
rect 26200 25072 26206 25084
rect 39850 25072 39856 25084
rect 26200 25044 39856 25072
rect 26200 25032 26206 25044
rect 39850 25032 39856 25044
rect 39908 25032 39914 25084
rect 9122 24964 9128 25016
rect 9180 25004 9186 25016
rect 17402 25004 17408 25016
rect 9180 24976 17408 25004
rect 9180 24964 9186 24976
rect 17402 24964 17408 24976
rect 17460 24964 17466 25016
rect 27154 24964 27160 25016
rect 27212 25004 27218 25016
rect 40034 25004 40040 25016
rect 27212 24976 40040 25004
rect 27212 24964 27218 24976
rect 40034 24964 40040 24976
rect 40092 24964 40098 25016
rect 28902 24896 28908 24948
rect 28960 24936 28966 24948
rect 35618 24936 35624 24948
rect 28960 24908 35624 24936
rect 28960 24896 28966 24908
rect 35618 24896 35624 24908
rect 35676 24896 35682 24948
rect 3142 24828 3148 24880
rect 3200 24868 3206 24880
rect 4430 24868 4436 24880
rect 3200 24840 4436 24868
rect 3200 24828 3206 24840
rect 4430 24828 4436 24840
rect 4488 24828 4494 24880
rect 7098 24828 7104 24880
rect 7156 24868 7162 24880
rect 15286 24868 15292 24880
rect 7156 24840 15292 24868
rect 7156 24828 7162 24840
rect 15286 24828 15292 24840
rect 15344 24868 15350 24880
rect 16666 24868 16672 24880
rect 15344 24840 16672 24868
rect 15344 24828 15350 24840
rect 16666 24828 16672 24840
rect 16724 24828 16730 24880
rect 28994 24828 29000 24880
rect 29052 24868 29058 24880
rect 40126 24868 40132 24880
rect 29052 24840 40132 24868
rect 29052 24828 29058 24840
rect 40126 24828 40132 24840
rect 40184 24828 40190 24880
rect 14274 24760 14280 24812
rect 14332 24800 14338 24812
rect 25498 24800 25504 24812
rect 14332 24772 25504 24800
rect 14332 24760 14338 24772
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 26602 24760 26608 24812
rect 26660 24800 26666 24812
rect 30098 24800 30104 24812
rect 26660 24772 30104 24800
rect 26660 24760 26666 24772
rect 30098 24760 30104 24772
rect 30156 24760 30162 24812
rect 35710 24760 35716 24812
rect 35768 24800 35774 24812
rect 38378 24800 38384 24812
rect 35768 24772 38384 24800
rect 35768 24760 35774 24772
rect 38378 24760 38384 24772
rect 38436 24760 38442 24812
rect 4338 24692 4344 24744
rect 4396 24732 4402 24744
rect 15010 24732 15016 24744
rect 4396 24704 15016 24732
rect 4396 24692 4402 24704
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 15378 24692 15384 24744
rect 15436 24732 15442 24744
rect 21174 24732 21180 24744
rect 15436 24704 21180 24732
rect 15436 24692 15442 24704
rect 21174 24692 21180 24704
rect 21232 24732 21238 24744
rect 27430 24732 27436 24744
rect 21232 24704 27436 24732
rect 21232 24692 21238 24704
rect 27430 24692 27436 24704
rect 27488 24692 27494 24744
rect 27522 24692 27528 24744
rect 27580 24732 27586 24744
rect 29086 24732 29092 24744
rect 27580 24704 29092 24732
rect 27580 24692 27586 24704
rect 29086 24692 29092 24704
rect 29144 24692 29150 24744
rect 31202 24692 31208 24744
rect 31260 24732 31266 24744
rect 37734 24732 37740 24744
rect 31260 24704 37740 24732
rect 31260 24692 31266 24704
rect 37734 24692 37740 24704
rect 37792 24692 37798 24744
rect 14918 24624 14924 24676
rect 14976 24664 14982 24676
rect 24486 24664 24492 24676
rect 14976 24636 24492 24664
rect 14976 24624 14982 24636
rect 24486 24624 24492 24636
rect 24544 24624 24550 24676
rect 29362 24664 29368 24676
rect 24780 24636 29368 24664
rect 3786 24556 3792 24608
rect 3844 24596 3850 24608
rect 21358 24596 21364 24608
rect 3844 24568 21364 24596
rect 3844 24556 3850 24568
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 24394 24556 24400 24608
rect 24452 24596 24458 24608
rect 24780 24596 24808 24636
rect 29362 24624 29368 24636
rect 29420 24624 29426 24676
rect 32214 24624 32220 24676
rect 32272 24664 32278 24676
rect 36630 24664 36636 24676
rect 32272 24636 36636 24664
rect 32272 24624 32278 24636
rect 36630 24624 36636 24636
rect 36688 24624 36694 24676
rect 24452 24568 24808 24596
rect 24452 24556 24458 24568
rect 24854 24556 24860 24608
rect 24912 24596 24918 24608
rect 27706 24596 27712 24608
rect 24912 24568 27712 24596
rect 24912 24556 24918 24568
rect 27706 24556 27712 24568
rect 27764 24556 27770 24608
rect 28074 24556 28080 24608
rect 28132 24596 28138 24608
rect 29178 24596 29184 24608
rect 28132 24568 29184 24596
rect 28132 24556 28138 24568
rect 29178 24556 29184 24568
rect 29236 24556 29242 24608
rect 29270 24556 29276 24608
rect 29328 24596 29334 24608
rect 36906 24596 36912 24608
rect 29328 24568 36912 24596
rect 29328 24556 29334 24568
rect 36906 24556 36912 24568
rect 36964 24556 36970 24608
rect 36998 24556 37004 24608
rect 37056 24596 37062 24608
rect 39298 24596 39304 24608
rect 37056 24568 39304 24596
rect 37056 24556 37062 24568
rect 39298 24556 39304 24568
rect 39356 24556 39362 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 3970 24352 3976 24404
rect 4028 24352 4034 24404
rect 4157 24395 4215 24401
rect 4157 24361 4169 24395
rect 4203 24392 4215 24395
rect 4246 24392 4252 24404
rect 4203 24364 4252 24392
rect 4203 24361 4215 24364
rect 4157 24355 4215 24361
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 4338 24352 4344 24404
rect 4396 24352 4402 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 24394 24392 24400 24404
rect 9171 24364 24400 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 24486 24352 24492 24404
rect 24544 24392 24550 24404
rect 24581 24395 24639 24401
rect 24581 24392 24593 24395
rect 24544 24364 24593 24392
rect 24544 24352 24550 24364
rect 24581 24361 24593 24364
rect 24627 24361 24639 24395
rect 24581 24355 24639 24361
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 31570 24392 31576 24404
rect 25188 24364 31576 24392
rect 25188 24352 25194 24364
rect 31570 24352 31576 24364
rect 31628 24352 31634 24404
rect 32858 24352 32864 24404
rect 32916 24392 32922 24404
rect 32953 24395 33011 24401
rect 32953 24392 32965 24395
rect 32916 24364 32965 24392
rect 32916 24352 32922 24364
rect 32953 24361 32965 24364
rect 32999 24361 33011 24395
rect 32953 24355 33011 24361
rect 35066 24352 35072 24404
rect 35124 24392 35130 24404
rect 38013 24395 38071 24401
rect 38013 24392 38025 24395
rect 35124 24364 38025 24392
rect 35124 24352 35130 24364
rect 38013 24361 38025 24364
rect 38059 24361 38071 24395
rect 38013 24355 38071 24361
rect 39298 24352 39304 24404
rect 39356 24352 39362 24404
rect 40034 24352 40040 24404
rect 40092 24352 40098 24404
rect 44726 24352 44732 24404
rect 44784 24352 44790 24404
rect 1578 24284 1584 24336
rect 1636 24284 1642 24336
rect 2774 24284 2780 24336
rect 2832 24324 2838 24336
rect 4706 24324 4712 24336
rect 2832 24296 4712 24324
rect 2832 24284 2838 24296
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 9306 24284 9312 24336
rect 9364 24284 9370 24336
rect 9398 24284 9404 24336
rect 9456 24324 9462 24336
rect 9456 24296 13492 24324
rect 9456 24284 9462 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 6822 24256 6828 24268
rect 5859 24228 6828 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9324 24256 9352 24284
rect 8251 24228 9352 24256
rect 10965 24259 11023 24265
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11011 24228 12434 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 1762 24148 1768 24200
rect 1820 24148 1826 24200
rect 2130 24148 2136 24200
rect 2188 24148 2194 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 2746 24160 4629 24188
rect 750 24080 756 24132
rect 808 24120 814 24132
rect 2746 24120 2774 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 9306 24148 9312 24200
rect 9364 24148 9370 24200
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10042 24188 10048 24200
rect 9999 24160 10048 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10042 24148 10048 24160
rect 10100 24148 10106 24200
rect 808 24092 2774 24120
rect 808 24080 814 24092
rect 3970 24080 3976 24132
rect 4028 24120 4034 24132
rect 7466 24120 7472 24132
rect 4028 24092 7472 24120
rect 4028 24080 4034 24092
rect 7466 24080 7472 24092
rect 7524 24080 7530 24132
rect 8938 24080 8944 24132
rect 8996 24120 9002 24132
rect 12406 24120 12434 24228
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 12618 24188 12624 24200
rect 12575 24160 12624 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 13464 24188 13492 24296
rect 14274 24284 14280 24336
rect 14332 24284 14338 24336
rect 18874 24284 18880 24336
rect 18932 24324 18938 24336
rect 18969 24327 19027 24333
rect 18969 24324 18981 24327
rect 18932 24296 18981 24324
rect 18932 24284 18938 24296
rect 18969 24293 18981 24296
rect 19015 24324 19027 24327
rect 23382 24324 23388 24336
rect 19015 24296 23388 24324
rect 19015 24293 19027 24296
rect 18969 24287 19027 24293
rect 23382 24284 23388 24296
rect 23440 24284 23446 24336
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 28905 24327 28963 24333
rect 28905 24324 28917 24327
rect 27672 24296 28917 24324
rect 27672 24284 27678 24296
rect 28905 24293 28917 24296
rect 28951 24293 28963 24327
rect 28905 24287 28963 24293
rect 29086 24284 29092 24336
rect 29144 24324 29150 24336
rect 29144 24296 30512 24324
rect 29144 24284 29150 24296
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 14366 24256 14372 24268
rect 13587 24228 14372 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 14366 24216 14372 24228
rect 14424 24216 14430 24268
rect 14734 24216 14740 24268
rect 14792 24256 14798 24268
rect 16853 24259 16911 24265
rect 14792 24228 16344 24256
rect 14792 24216 14798 24228
rect 13464 24160 14412 24188
rect 13814 24120 13820 24132
rect 8996 24092 11928 24120
rect 12406 24092 13820 24120
rect 8996 24080 9002 24092
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 9490 24052 9496 24064
rect 6595 24024 9496 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 9490 24012 9496 24024
rect 9548 24012 9554 24064
rect 11698 24012 11704 24064
rect 11756 24052 11762 24064
rect 11793 24055 11851 24061
rect 11793 24052 11805 24055
rect 11756 24024 11805 24052
rect 11756 24012 11762 24024
rect 11793 24021 11805 24024
rect 11839 24021 11851 24055
rect 11900 24052 11928 24092
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 14384 24120 14412 24160
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 14826 24148 14832 24200
rect 14884 24188 14890 24200
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14884 24160 14933 24188
rect 14884 24148 14890 24160
rect 14921 24157 14933 24160
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 16022 24120 16028 24132
rect 14384 24092 16028 24120
rect 16022 24080 16028 24092
rect 16080 24080 16086 24132
rect 16117 24123 16175 24129
rect 16117 24089 16129 24123
rect 16163 24120 16175 24123
rect 16206 24120 16212 24132
rect 16163 24092 16212 24120
rect 16163 24089 16175 24092
rect 16117 24083 16175 24089
rect 16206 24080 16212 24092
rect 16264 24080 16270 24132
rect 16316 24120 16344 24228
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 17126 24256 17132 24268
rect 16899 24228 17132 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21600 24228 22477 24256
rect 21600 24216 21606 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 25038 24256 25044 24268
rect 22465 24219 22523 24225
rect 24872 24228 25044 24256
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 24872 24188 24900 24228
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 25222 24216 25228 24268
rect 25280 24216 25286 24268
rect 26326 24216 26332 24268
rect 26384 24216 26390 24268
rect 26970 24216 26976 24268
rect 27028 24256 27034 24268
rect 28074 24256 28080 24268
rect 27028 24228 28080 24256
rect 27028 24216 27034 24228
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 28350 24216 28356 24268
rect 28408 24216 28414 24268
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29733 24259 29791 24265
rect 29733 24256 29745 24259
rect 29328 24228 29745 24256
rect 29328 24216 29334 24228
rect 29733 24225 29745 24228
rect 29779 24225 29791 24259
rect 30484 24256 30512 24296
rect 30558 24284 30564 24336
rect 30616 24324 30622 24336
rect 30616 24296 40264 24324
rect 30616 24284 30622 24296
rect 31662 24256 31668 24268
rect 30484 24228 31668 24256
rect 29733 24219 29791 24225
rect 31662 24216 31668 24228
rect 31720 24216 31726 24268
rect 33042 24216 33048 24268
rect 33100 24256 33106 24268
rect 35529 24259 35587 24265
rect 35529 24256 35541 24259
rect 33100 24228 35541 24256
rect 33100 24216 33106 24228
rect 35529 24225 35541 24228
rect 35575 24225 35587 24259
rect 35529 24219 35587 24225
rect 35728 24228 38608 24256
rect 22235 24160 24900 24188
rect 24949 24191 25007 24197
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 24949 24157 24961 24191
rect 24995 24188 25007 24191
rect 25314 24188 25320 24200
rect 24995 24160 25320 24188
rect 24995 24157 25007 24160
rect 24949 24151 25007 24157
rect 25314 24148 25320 24160
rect 25372 24148 25378 24200
rect 26142 24148 26148 24200
rect 26200 24188 26206 24200
rect 26237 24191 26295 24197
rect 26237 24188 26249 24191
rect 26200 24160 26249 24188
rect 26200 24148 26206 24160
rect 26237 24157 26249 24160
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 26418 24148 26424 24200
rect 26476 24188 26482 24200
rect 26476 24160 28672 24188
rect 26476 24148 26482 24160
rect 17129 24123 17187 24129
rect 17129 24120 17141 24123
rect 16316 24092 17141 24120
rect 17129 24089 17141 24092
rect 17175 24089 17187 24123
rect 18414 24120 18420 24132
rect 18354 24092 18420 24120
rect 17129 24083 17187 24089
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 19518 24080 19524 24132
rect 19576 24120 19582 24132
rect 19576 24092 25820 24120
rect 19576 24080 19582 24092
rect 11977 24055 12035 24061
rect 11977 24052 11989 24055
rect 11900 24024 11989 24052
rect 11793 24015 11851 24021
rect 11977 24021 11989 24024
rect 12023 24052 12035 24055
rect 15378 24052 15384 24064
rect 12023 24024 15384 24052
rect 12023 24021 12035 24024
rect 11977 24015 12035 24021
rect 15378 24012 15384 24024
rect 15436 24012 15442 24064
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 15528 24024 18613 24052
rect 15528 24012 15534 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 23658 24052 23664 24064
rect 19475 24024 23664 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24052 23903 24055
rect 24762 24052 24768 24064
rect 23891 24024 24768 24052
rect 23891 24021 23903 24024
rect 23845 24015 23903 24021
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25682 24052 25688 24064
rect 25087 24024 25688 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25682 24012 25688 24024
rect 25740 24012 25746 24064
rect 25792 24061 25820 24092
rect 26786 24080 26792 24132
rect 26844 24120 26850 24132
rect 27341 24123 27399 24129
rect 27341 24120 27353 24123
rect 26844 24092 27353 24120
rect 26844 24080 26850 24092
rect 27341 24089 27353 24092
rect 27387 24120 27399 24123
rect 27798 24120 27804 24132
rect 27387 24092 27804 24120
rect 27387 24089 27399 24092
rect 27341 24083 27399 24089
rect 27798 24080 27804 24092
rect 27856 24120 27862 24132
rect 28534 24120 28540 24132
rect 27856 24092 28540 24120
rect 27856 24080 27862 24092
rect 28534 24080 28540 24092
rect 28592 24080 28598 24132
rect 28644 24120 28672 24160
rect 29086 24148 29092 24200
rect 29144 24148 29150 24200
rect 29822 24148 29828 24200
rect 29880 24188 29886 24200
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 29880 24160 30021 24188
rect 29880 24148 29886 24160
rect 30009 24157 30021 24160
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 30098 24148 30104 24200
rect 30156 24188 30162 24200
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 30156 24160 31033 24188
rect 30156 24148 30162 24160
rect 31021 24157 31033 24160
rect 31067 24157 31079 24191
rect 31021 24151 31079 24157
rect 31110 24148 31116 24200
rect 31168 24188 31174 24200
rect 32309 24191 32367 24197
rect 32309 24188 32321 24191
rect 31168 24160 32321 24188
rect 31168 24148 31174 24160
rect 32309 24157 32321 24160
rect 32355 24157 32367 24191
rect 32309 24151 32367 24157
rect 33413 24191 33471 24197
rect 33413 24157 33425 24191
rect 33459 24157 33471 24191
rect 33413 24151 33471 24157
rect 33428 24120 33456 24151
rect 33870 24148 33876 24200
rect 33928 24188 33934 24200
rect 34333 24191 34391 24197
rect 34333 24188 34345 24191
rect 33928 24160 34345 24188
rect 33928 24148 33934 24160
rect 34333 24157 34345 24160
rect 34379 24157 34391 24191
rect 34333 24151 34391 24157
rect 34882 24148 34888 24200
rect 34940 24188 34946 24200
rect 35728 24188 35756 24228
rect 34940 24160 35756 24188
rect 34940 24148 34946 24160
rect 35802 24148 35808 24200
rect 35860 24188 35866 24200
rect 36909 24191 36967 24197
rect 36909 24188 36921 24191
rect 35860 24160 36921 24188
rect 35860 24148 35866 24160
rect 36909 24157 36921 24160
rect 36955 24188 36967 24191
rect 36955 24160 37688 24188
rect 36955 24157 36967 24160
rect 36909 24151 36967 24157
rect 28644 24092 33456 24120
rect 33502 24080 33508 24132
rect 33560 24120 33566 24132
rect 36081 24123 36139 24129
rect 36081 24120 36093 24123
rect 33560 24092 36093 24120
rect 33560 24080 33566 24092
rect 35820 24064 35848 24092
rect 36081 24089 36093 24092
rect 36127 24089 36139 24123
rect 36081 24083 36139 24089
rect 37366 24080 37372 24132
rect 37424 24120 37430 24132
rect 37553 24123 37611 24129
rect 37553 24120 37565 24123
rect 37424 24092 37565 24120
rect 37424 24080 37430 24092
rect 37553 24089 37565 24092
rect 37599 24089 37611 24123
rect 37660 24120 37688 24160
rect 38286 24148 38292 24200
rect 38344 24188 38350 24200
rect 38473 24191 38531 24197
rect 38473 24188 38485 24191
rect 38344 24160 38485 24188
rect 38344 24148 38350 24160
rect 38473 24157 38485 24160
rect 38519 24157 38531 24191
rect 38473 24151 38531 24157
rect 38580 24120 38608 24228
rect 38654 24216 38660 24268
rect 38712 24216 38718 24268
rect 40236 24256 40264 24296
rect 43530 24284 43536 24336
rect 43588 24324 43594 24336
rect 46845 24327 46903 24333
rect 46845 24324 46857 24327
rect 43588 24296 46857 24324
rect 43588 24284 43594 24296
rect 46845 24293 46857 24296
rect 46891 24293 46903 24327
rect 46845 24287 46903 24293
rect 40236 24228 41414 24256
rect 38930 24148 38936 24200
rect 38988 24188 38994 24200
rect 39206 24188 39212 24200
rect 38988 24160 39212 24188
rect 38988 24148 38994 24160
rect 39206 24148 39212 24160
rect 39264 24148 39270 24200
rect 40236 24197 40264 24228
rect 40221 24191 40279 24197
rect 40221 24157 40233 24191
rect 40267 24157 40279 24191
rect 40221 24151 40279 24157
rect 40310 24148 40316 24200
rect 40368 24188 40374 24200
rect 41230 24188 41236 24200
rect 40368 24160 41236 24188
rect 40368 24148 40374 24160
rect 41230 24148 41236 24160
rect 41288 24148 41294 24200
rect 41386 24188 41414 24228
rect 41386 24160 41460 24188
rect 40497 24123 40555 24129
rect 40497 24120 40509 24123
rect 37660 24092 38148 24120
rect 38580 24092 40509 24120
rect 37553 24083 37611 24089
rect 25777 24055 25835 24061
rect 25777 24021 25789 24055
rect 25823 24021 25835 24055
rect 25777 24015 25835 24021
rect 25958 24012 25964 24064
rect 26016 24052 26022 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 26016 24024 26157 24052
rect 26016 24012 26022 24024
rect 26145 24021 26157 24024
rect 26191 24052 26203 24055
rect 26970 24052 26976 24064
rect 26191 24024 26976 24052
rect 26191 24021 26203 24024
rect 26145 24015 26203 24021
rect 26970 24012 26976 24024
rect 27028 24012 27034 24064
rect 27246 24012 27252 24064
rect 27304 24012 27310 24064
rect 27706 24012 27712 24064
rect 27764 24012 27770 24064
rect 28074 24012 28080 24064
rect 28132 24012 28138 24064
rect 28169 24055 28227 24061
rect 28169 24021 28181 24055
rect 28215 24052 28227 24055
rect 28810 24052 28816 24064
rect 28215 24024 28816 24052
rect 28215 24021 28227 24024
rect 28169 24015 28227 24021
rect 28810 24012 28816 24024
rect 28868 24012 28874 24064
rect 28994 24012 29000 24064
rect 29052 24052 29058 24064
rect 31665 24055 31723 24061
rect 31665 24052 31677 24055
rect 29052 24024 31677 24052
rect 29052 24012 29058 24024
rect 31665 24021 31677 24024
rect 31711 24021 31723 24055
rect 31665 24015 31723 24021
rect 32766 24012 32772 24064
rect 32824 24052 32830 24064
rect 34057 24055 34115 24061
rect 34057 24052 34069 24055
rect 32824 24024 34069 24052
rect 32824 24012 32830 24024
rect 34057 24021 34069 24024
rect 34103 24021 34115 24055
rect 34057 24015 34115 24021
rect 35802 24012 35808 24064
rect 35860 24012 35866 24064
rect 35986 24012 35992 24064
rect 36044 24052 36050 24064
rect 36173 24055 36231 24061
rect 36173 24052 36185 24055
rect 36044 24024 36185 24052
rect 36044 24012 36050 24024
rect 36173 24021 36185 24024
rect 36219 24021 36231 24055
rect 36173 24015 36231 24021
rect 36722 24012 36728 24064
rect 36780 24012 36786 24064
rect 37274 24012 37280 24064
rect 37332 24052 37338 24064
rect 37645 24055 37703 24061
rect 37645 24052 37657 24055
rect 37332 24024 37657 24052
rect 37332 24012 37338 24024
rect 37645 24021 37657 24024
rect 37691 24021 37703 24055
rect 38120 24052 38148 24092
rect 40497 24089 40509 24092
rect 40543 24089 40555 24123
rect 41432 24120 41460 24160
rect 41506 24148 41512 24200
rect 41564 24148 41570 24200
rect 41598 24148 41604 24200
rect 41656 24188 41662 24200
rect 42610 24188 42616 24200
rect 41656 24160 42616 24188
rect 41656 24148 41662 24160
rect 42610 24148 42616 24160
rect 42668 24148 42674 24200
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44784 24160 45201 24188
rect 44784 24148 44790 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24157 45983 24191
rect 45925 24151 45983 24157
rect 46014 24148 46020 24200
rect 46072 24188 46078 24200
rect 46661 24191 46719 24197
rect 46661 24188 46673 24191
rect 46072 24160 46673 24188
rect 46072 24148 46078 24160
rect 46661 24157 46673 24160
rect 46707 24188 46719 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 46707 24160 47225 24188
rect 46707 24157 46719 24160
rect 46661 24151 46719 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 47946 24148 47952 24200
rect 48004 24188 48010 24200
rect 48501 24191 48559 24197
rect 48501 24188 48513 24191
rect 48004 24160 48513 24188
rect 48004 24148 48010 24160
rect 48501 24157 48513 24160
rect 48547 24188 48559 24191
rect 49053 24191 49111 24197
rect 49053 24188 49065 24191
rect 48547 24160 49065 24188
rect 48547 24157 48559 24160
rect 48501 24151 48559 24157
rect 49053 24157 49065 24160
rect 49099 24157 49111 24191
rect 49053 24151 49111 24157
rect 42426 24120 42432 24132
rect 41432 24092 42432 24120
rect 40497 24083 40555 24089
rect 42426 24080 42432 24092
rect 42484 24080 42490 24132
rect 42518 24080 42524 24132
rect 42576 24120 42582 24132
rect 42576 24092 45554 24120
rect 42576 24080 42582 24092
rect 40681 24055 40739 24061
rect 40681 24052 40693 24055
rect 38120 24024 40693 24052
rect 37645 24015 37703 24021
rect 40681 24021 40693 24024
rect 40727 24021 40739 24055
rect 40681 24015 40739 24021
rect 40770 24012 40776 24064
rect 40828 24052 40834 24064
rect 40865 24055 40923 24061
rect 40865 24052 40877 24055
rect 40828 24024 40877 24052
rect 40828 24012 40834 24024
rect 40865 24021 40877 24024
rect 40911 24021 40923 24055
rect 40865 24015 40923 24021
rect 43898 24012 43904 24064
rect 43956 24012 43962 24064
rect 45278 24012 45284 24064
rect 45336 24052 45342 24064
rect 45373 24055 45431 24061
rect 45373 24052 45385 24055
rect 45336 24024 45385 24052
rect 45336 24012 45342 24024
rect 45373 24021 45385 24024
rect 45419 24021 45431 24055
rect 45526 24052 45554 24092
rect 46109 24055 46167 24061
rect 46109 24052 46121 24055
rect 45526 24024 46121 24052
rect 45373 24015 45431 24021
rect 46109 24021 46121 24024
rect 46155 24021 46167 24055
rect 46109 24015 46167 24021
rect 47026 24012 47032 24064
rect 47084 24052 47090 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 47084 24024 47961 24052
rect 47084 24012 47090 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 48590 24012 48596 24064
rect 48648 24052 48654 24064
rect 48685 24055 48743 24061
rect 48685 24052 48697 24055
rect 48648 24024 48697 24052
rect 48648 24012 48654 24024
rect 48685 24021 48697 24024
rect 48731 24021 48743 24055
rect 48685 24015 48743 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 9398 23848 9404 23860
rect 2148 23820 9404 23848
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 2148 23712 2176 23820
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 15470 23848 15476 23860
rect 10192 23820 15476 23848
rect 10192 23808 10198 23820
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 16761 23851 16819 23857
rect 16761 23817 16773 23851
rect 16807 23848 16819 23851
rect 22278 23848 22284 23860
rect 16807 23820 22284 23848
rect 16807 23817 16819 23820
rect 16761 23811 16819 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22646 23808 22652 23860
rect 22704 23848 22710 23860
rect 26970 23848 26976 23860
rect 22704 23820 26976 23848
rect 22704 23808 22710 23820
rect 26970 23808 26976 23820
rect 27028 23808 27034 23860
rect 27080 23820 28764 23848
rect 2406 23740 2412 23792
rect 2464 23780 2470 23792
rect 7101 23783 7159 23789
rect 2464 23752 4660 23780
rect 2464 23740 2470 23752
rect 1719 23684 2176 23712
rect 2777 23715 2835 23721
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2777 23681 2789 23715
rect 2823 23681 2835 23715
rect 2777 23675 2835 23681
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23712 4031 23715
rect 4154 23712 4160 23724
rect 4019 23684 4160 23712
rect 4019 23681 4031 23684
rect 3973 23675 4031 23681
rect 842 23604 848 23656
rect 900 23644 906 23656
rect 2792 23644 2820 23675
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4632 23721 4660 23752
rect 7101 23749 7113 23783
rect 7147 23780 7159 23783
rect 9125 23783 9183 23789
rect 7147 23752 8708 23780
rect 7147 23749 7159 23752
rect 7101 23743 7159 23749
rect 4617 23715 4675 23721
rect 4617 23681 4629 23715
rect 4663 23681 4675 23715
rect 4617 23675 4675 23681
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23712 7251 23715
rect 7650 23712 7656 23724
rect 7239 23684 7656 23712
rect 7239 23681 7251 23684
rect 7193 23675 7251 23681
rect 7650 23672 7656 23684
rect 7708 23672 7714 23724
rect 8110 23672 8116 23724
rect 8168 23672 8174 23724
rect 900 23616 2820 23644
rect 900 23604 906 23616
rect 3694 23604 3700 23656
rect 3752 23644 3758 23656
rect 4522 23644 4528 23656
rect 3752 23616 4528 23644
rect 3752 23604 3758 23616
rect 4522 23604 4528 23616
rect 4580 23604 4586 23656
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23644 7435 23647
rect 7558 23644 7564 23656
rect 7423 23616 7564 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 8680 23644 8708 23752
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9950 23780 9956 23792
rect 9171 23752 9956 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 12526 23780 12532 23792
rect 11011 23752 12532 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 12526 23740 12532 23752
rect 12584 23740 12590 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23780 18291 23783
rect 19058 23780 19064 23792
rect 18279 23752 19064 23780
rect 18279 23749 18291 23752
rect 18233 23743 18291 23749
rect 19058 23740 19064 23752
rect 19116 23740 19122 23792
rect 19153 23783 19211 23789
rect 19153 23749 19165 23783
rect 19199 23780 19211 23783
rect 19242 23780 19248 23792
rect 19199 23752 19248 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 20438 23780 20444 23792
rect 20378 23752 20444 23780
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 21358 23740 21364 23792
rect 21416 23740 21422 23792
rect 23566 23780 23572 23792
rect 23506 23752 23572 23780
rect 23566 23740 23572 23752
rect 23624 23740 23630 23792
rect 25130 23740 25136 23792
rect 25188 23740 25194 23792
rect 26786 23780 26792 23792
rect 26358 23752 26792 23780
rect 26786 23740 26792 23752
rect 26844 23740 26850 23792
rect 9858 23672 9864 23724
rect 9916 23672 9922 23724
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23712 11759 23715
rect 13265 23715 13323 23721
rect 11747 23684 12434 23712
rect 11747 23681 11759 23684
rect 11701 23675 11759 23681
rect 10226 23644 10232 23656
rect 8680 23616 10232 23644
rect 10226 23604 10232 23616
rect 10284 23604 10290 23656
rect 11974 23604 11980 23656
rect 12032 23604 12038 23656
rect 12406 23644 12434 23684
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13722 23712 13728 23724
rect 13311 23684 13728 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 14734 23712 14740 23724
rect 14568 23684 14740 23712
rect 14366 23644 14372 23656
rect 12406 23616 14372 23644
rect 14366 23604 14372 23616
rect 14424 23604 14430 23656
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 14568 23576 14596 23684
rect 14734 23672 14740 23684
rect 14792 23672 14798 23724
rect 15010 23672 15016 23724
rect 15068 23672 15074 23724
rect 16942 23712 16948 23724
rect 15948 23684 16948 23712
rect 15948 23644 15976 23684
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 17221 23715 17279 23721
rect 17221 23681 17233 23715
rect 17267 23712 17279 23715
rect 17402 23712 17408 23724
rect 17267 23684 17408 23712
rect 17267 23681 17279 23684
rect 17221 23675 17279 23681
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 21174 23672 21180 23724
rect 21232 23672 21238 23724
rect 2363 23548 14596 23576
rect 14660 23616 15976 23644
rect 16117 23647 16175 23653
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 566 23468 572 23520
rect 624 23508 630 23520
rect 2406 23508 2412 23520
rect 624 23480 2412 23508
rect 624 23468 630 23480
rect 2406 23468 2412 23480
rect 2464 23468 2470 23520
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 6365 23511 6423 23517
rect 6365 23508 6377 23511
rect 5592 23480 6377 23508
rect 5592 23468 5598 23480
rect 6365 23477 6377 23480
rect 6411 23508 6423 23511
rect 6546 23508 6552 23520
rect 6411 23480 6552 23508
rect 6411 23477 6423 23480
rect 6365 23471 6423 23477
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 6733 23511 6791 23517
rect 6733 23508 6745 23511
rect 6696 23480 6745 23508
rect 6696 23468 6702 23480
rect 6733 23477 6745 23480
rect 6779 23477 6791 23511
rect 6733 23471 6791 23477
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 14660 23508 14688 23616
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 16298 23644 16304 23656
rect 16163 23616 16304 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 16298 23604 16304 23616
rect 16356 23604 16362 23656
rect 18877 23647 18935 23653
rect 18877 23613 18889 23647
rect 18923 23644 18935 23647
rect 18923 23616 19012 23644
rect 18923 23613 18935 23616
rect 18877 23607 18935 23613
rect 9548 23480 14688 23508
rect 18984 23508 19012 23616
rect 20346 23604 20352 23656
rect 20404 23644 20410 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20404 23616 22017 23644
rect 20404 23604 20410 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22281 23647 22339 23653
rect 22281 23613 22293 23647
rect 22327 23644 22339 23647
rect 22646 23644 22652 23656
rect 22327 23616 22652 23644
rect 22327 23613 22339 23616
rect 22281 23607 22339 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 22830 23604 22836 23656
rect 22888 23644 22894 23656
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 22888 23616 24225 23644
rect 22888 23604 22894 23616
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 24857 23647 24915 23653
rect 24857 23613 24869 23647
rect 24903 23613 24915 23647
rect 24857 23607 24915 23613
rect 23290 23536 23296 23588
rect 23348 23576 23354 23588
rect 24872 23576 24900 23607
rect 25682 23604 25688 23656
rect 25740 23644 25746 23656
rect 27080 23644 27108 23820
rect 27430 23740 27436 23792
rect 27488 23780 27494 23792
rect 27706 23780 27712 23792
rect 27488 23752 27712 23780
rect 27488 23740 27494 23752
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 27890 23740 27896 23792
rect 27948 23740 27954 23792
rect 28736 23780 28764 23820
rect 28810 23808 28816 23860
rect 28868 23848 28874 23860
rect 28868 23820 32812 23848
rect 28868 23808 28874 23820
rect 30190 23780 30196 23792
rect 28736 23752 30196 23780
rect 30190 23740 30196 23752
rect 30248 23740 30254 23792
rect 30374 23740 30380 23792
rect 30432 23780 30438 23792
rect 30742 23780 30748 23792
rect 30432 23752 30748 23780
rect 30432 23740 30438 23752
rect 30742 23740 30748 23752
rect 30800 23740 30806 23792
rect 32784 23780 32812 23820
rect 32858 23808 32864 23860
rect 32916 23848 32922 23860
rect 33965 23851 34023 23857
rect 33965 23848 33977 23851
rect 32916 23820 33977 23848
rect 32916 23808 32922 23820
rect 33965 23817 33977 23820
rect 34011 23817 34023 23851
rect 33965 23811 34023 23817
rect 36538 23808 36544 23860
rect 36596 23808 36602 23860
rect 36906 23808 36912 23860
rect 36964 23808 36970 23860
rect 37458 23808 37464 23860
rect 37516 23808 37522 23860
rect 38746 23808 38752 23860
rect 38804 23848 38810 23860
rect 38933 23851 38991 23857
rect 38933 23848 38945 23851
rect 38804 23820 38945 23848
rect 38804 23808 38810 23820
rect 38933 23817 38945 23820
rect 38979 23817 38991 23851
rect 38933 23811 38991 23817
rect 39206 23808 39212 23860
rect 39264 23848 39270 23860
rect 42153 23851 42211 23857
rect 42153 23848 42165 23851
rect 39264 23820 42165 23848
rect 39264 23808 39270 23820
rect 42153 23817 42165 23820
rect 42199 23817 42211 23851
rect 42153 23811 42211 23817
rect 42426 23808 42432 23860
rect 42484 23808 42490 23860
rect 42610 23808 42616 23860
rect 42668 23848 42674 23860
rect 42981 23851 43039 23857
rect 42981 23848 42993 23851
rect 42668 23820 42993 23848
rect 42668 23808 42674 23820
rect 42981 23817 42993 23820
rect 43027 23817 43039 23851
rect 42981 23811 43039 23817
rect 43257 23851 43315 23857
rect 43257 23817 43269 23851
rect 43303 23848 43315 23851
rect 43438 23848 43444 23860
rect 43303 23820 43444 23848
rect 43303 23817 43315 23820
rect 43257 23811 43315 23817
rect 43438 23808 43444 23820
rect 43496 23848 43502 23860
rect 43496 23820 43668 23848
rect 43496 23808 43502 23820
rect 40770 23780 40776 23792
rect 30852 23752 32352 23780
rect 32784 23752 36952 23780
rect 28718 23672 28724 23724
rect 28776 23712 28782 23724
rect 29641 23715 29699 23721
rect 29641 23712 29653 23715
rect 28776 23684 29653 23712
rect 28776 23672 28782 23684
rect 29641 23681 29653 23684
rect 29687 23681 29699 23715
rect 29641 23675 29699 23681
rect 30098 23672 30104 23724
rect 30156 23712 30162 23724
rect 30852 23712 30880 23752
rect 30156 23684 30880 23712
rect 30156 23672 30162 23684
rect 30926 23672 30932 23724
rect 30984 23672 30990 23724
rect 31018 23672 31024 23724
rect 31076 23712 31082 23724
rect 31573 23715 31631 23721
rect 31573 23712 31585 23715
rect 31076 23684 31585 23712
rect 31076 23672 31082 23684
rect 31573 23681 31585 23684
rect 31619 23712 31631 23715
rect 32214 23712 32220 23724
rect 31619 23684 32220 23712
rect 31619 23681 31631 23684
rect 31573 23675 31631 23681
rect 32214 23672 32220 23684
rect 32272 23672 32278 23724
rect 32324 23721 32352 23752
rect 36924 23724 36952 23752
rect 38304 23752 40776 23780
rect 32320 23715 32378 23721
rect 32320 23681 32332 23715
rect 32366 23681 32378 23715
rect 32320 23675 32378 23681
rect 34606 23672 34612 23724
rect 34664 23672 34670 23724
rect 35710 23721 35716 23724
rect 35696 23716 35716 23721
rect 35636 23715 35716 23716
rect 35636 23684 35708 23715
rect 25740 23616 27108 23644
rect 27157 23647 27215 23653
rect 25740 23604 25746 23616
rect 27157 23613 27169 23647
rect 27203 23613 27215 23647
rect 27157 23607 27215 23613
rect 27433 23647 27491 23653
rect 27433 23613 27445 23647
rect 27479 23644 27491 23647
rect 28994 23644 29000 23656
rect 27479 23616 29000 23644
rect 27479 23613 27491 23616
rect 27433 23607 27491 23613
rect 23348 23548 24900 23576
rect 23348 23536 23354 23548
rect 26602 23536 26608 23588
rect 26660 23536 26666 23588
rect 19702 23508 19708 23520
rect 18984 23480 19708 23508
rect 9548 23468 9554 23480
rect 19702 23468 19708 23480
rect 19760 23468 19766 23520
rect 19794 23468 19800 23520
rect 19852 23508 19858 23520
rect 20625 23511 20683 23517
rect 20625 23508 20637 23511
rect 19852 23480 20637 23508
rect 19852 23468 19858 23480
rect 20625 23477 20637 23480
rect 20671 23477 20683 23511
rect 20625 23471 20683 23477
rect 23753 23511 23811 23517
rect 23753 23477 23765 23511
rect 23799 23508 23811 23511
rect 26418 23508 26424 23520
rect 23799 23480 26424 23508
rect 23799 23477 23811 23480
rect 23753 23471 23811 23477
rect 26418 23468 26424 23480
rect 26476 23468 26482 23520
rect 27172 23508 27200 23607
rect 28994 23604 29000 23616
rect 29052 23604 29058 23656
rect 29362 23604 29368 23656
rect 29420 23604 29426 23656
rect 30006 23604 30012 23656
rect 30064 23644 30070 23656
rect 32953 23647 33011 23653
rect 32953 23644 32965 23647
rect 30064 23616 32965 23644
rect 30064 23604 30070 23616
rect 32953 23613 32965 23616
rect 32999 23613 33011 23647
rect 32953 23607 33011 23613
rect 34330 23604 34336 23656
rect 34388 23604 34394 23656
rect 34422 23604 34428 23656
rect 34480 23644 34486 23656
rect 35636 23644 35664 23684
rect 35696 23681 35708 23684
rect 35696 23675 35716 23681
rect 35710 23672 35716 23675
rect 35768 23672 35774 23724
rect 35894 23672 35900 23724
rect 35952 23672 35958 23724
rect 36446 23672 36452 23724
rect 36504 23672 36510 23724
rect 36906 23672 36912 23724
rect 36964 23672 36970 23724
rect 37734 23672 37740 23724
rect 37792 23712 37798 23724
rect 38304 23721 38332 23752
rect 40770 23740 40776 23752
rect 40828 23740 40834 23792
rect 41230 23740 41236 23792
rect 41288 23780 41294 23792
rect 43640 23789 43668 23820
rect 45554 23808 45560 23860
rect 45612 23848 45618 23860
rect 45741 23851 45799 23857
rect 45741 23848 45753 23851
rect 45612 23820 45753 23848
rect 45612 23808 45618 23820
rect 45741 23817 45753 23820
rect 45787 23817 45799 23851
rect 45741 23811 45799 23817
rect 47302 23808 47308 23860
rect 47360 23848 47366 23860
rect 47581 23851 47639 23857
rect 47581 23848 47593 23851
rect 47360 23820 47593 23848
rect 47360 23808 47366 23820
rect 47581 23817 47593 23820
rect 47627 23817 47639 23851
rect 47581 23811 47639 23817
rect 42797 23783 42855 23789
rect 42797 23780 42809 23783
rect 41288 23752 42809 23780
rect 41288 23740 41294 23752
rect 42797 23749 42809 23752
rect 42843 23749 42855 23783
rect 42797 23743 42855 23749
rect 43625 23783 43683 23789
rect 43625 23749 43637 23783
rect 43671 23749 43683 23783
rect 43625 23743 43683 23749
rect 38289 23715 38347 23721
rect 38289 23712 38301 23715
rect 37792 23684 38301 23712
rect 37792 23672 37798 23684
rect 38289 23681 38301 23684
rect 38335 23681 38347 23715
rect 38289 23675 38347 23681
rect 38841 23715 38899 23721
rect 38841 23681 38853 23715
rect 38887 23712 38899 23715
rect 39206 23712 39212 23724
rect 38887 23684 39212 23712
rect 38887 23681 38899 23684
rect 38841 23675 38899 23681
rect 39206 23672 39212 23684
rect 39264 23712 39270 23724
rect 39942 23712 39948 23724
rect 39264 23684 39948 23712
rect 39264 23672 39270 23684
rect 39942 23672 39948 23684
rect 40000 23672 40006 23724
rect 40037 23715 40095 23721
rect 40037 23681 40049 23715
rect 40083 23712 40095 23715
rect 40126 23712 40132 23724
rect 40083 23684 40132 23712
rect 40083 23681 40095 23684
rect 40037 23675 40095 23681
rect 40126 23672 40132 23684
rect 40184 23672 40190 23724
rect 40221 23715 40279 23721
rect 40221 23681 40233 23715
rect 40267 23712 40279 23715
rect 40402 23712 40408 23724
rect 40267 23684 40408 23712
rect 40267 23681 40279 23684
rect 40221 23675 40279 23681
rect 40402 23672 40408 23684
rect 40460 23672 40466 23724
rect 42613 23715 42671 23721
rect 42613 23712 42625 23715
rect 40696 23684 42625 23712
rect 34480 23616 35664 23644
rect 34480 23604 34486 23616
rect 35802 23604 35808 23656
rect 35860 23644 35866 23656
rect 39485 23647 39543 23653
rect 39485 23644 39497 23647
rect 35860 23616 39497 23644
rect 35860 23604 35866 23616
rect 39485 23613 39497 23616
rect 39531 23613 39543 23647
rect 39485 23607 39543 23613
rect 39574 23604 39580 23656
rect 39632 23644 39638 23656
rect 40696 23653 40724 23684
rect 42613 23681 42625 23684
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 44174 23672 44180 23724
rect 44232 23712 44238 23724
rect 44269 23715 44327 23721
rect 44269 23712 44281 23715
rect 44232 23684 44281 23712
rect 44232 23672 44238 23684
rect 44269 23681 44281 23684
rect 44315 23712 44327 23715
rect 44821 23715 44879 23721
rect 44821 23712 44833 23715
rect 44315 23684 44833 23712
rect 44315 23681 44327 23684
rect 44269 23675 44327 23681
rect 44821 23681 44833 23684
rect 44867 23681 44879 23715
rect 44821 23675 44879 23681
rect 46658 23672 46664 23724
rect 46716 23712 46722 23724
rect 46753 23715 46811 23721
rect 46753 23712 46765 23715
rect 46716 23684 46765 23712
rect 46716 23672 46722 23684
rect 46753 23681 46765 23684
rect 46799 23712 46811 23715
rect 47305 23715 47363 23721
rect 47305 23712 47317 23715
rect 46799 23684 47317 23712
rect 46799 23681 46811 23684
rect 46753 23675 46811 23681
rect 47305 23681 47317 23684
rect 47351 23681 47363 23715
rect 47305 23675 47363 23681
rect 48866 23672 48872 23724
rect 48924 23712 48930 23724
rect 49145 23715 49203 23721
rect 49145 23712 49157 23715
rect 48924 23684 49157 23712
rect 48924 23672 48930 23684
rect 49145 23681 49157 23684
rect 49191 23681 49203 23715
rect 49145 23675 49203 23681
rect 40681 23647 40739 23653
rect 40681 23644 40693 23647
rect 39632 23616 40693 23644
rect 39632 23604 39638 23616
rect 40681 23613 40693 23616
rect 40727 23613 40739 23647
rect 40681 23607 40739 23613
rect 40954 23604 40960 23656
rect 41012 23604 41018 23656
rect 41046 23604 41052 23656
rect 41104 23644 41110 23656
rect 41969 23647 42027 23653
rect 41969 23644 41981 23647
rect 41104 23616 41981 23644
rect 41104 23604 41110 23616
rect 41969 23613 41981 23616
rect 42015 23613 42027 23647
rect 41969 23607 42027 23613
rect 29270 23576 29276 23588
rect 28460 23548 29276 23576
rect 27522 23508 27528 23520
rect 27172 23480 27528 23508
rect 27522 23468 27528 23480
rect 27580 23468 27586 23520
rect 27798 23468 27804 23520
rect 27856 23508 27862 23520
rect 28460 23508 28488 23548
rect 29270 23536 29276 23548
rect 29328 23536 29334 23588
rect 31662 23536 31668 23588
rect 31720 23576 31726 23588
rect 33413 23579 33471 23585
rect 33413 23576 33425 23579
rect 31720 23548 33425 23576
rect 31720 23536 31726 23548
rect 33413 23545 33425 23548
rect 33459 23545 33471 23579
rect 33413 23539 33471 23545
rect 33689 23579 33747 23585
rect 33689 23545 33701 23579
rect 33735 23576 33747 23579
rect 33870 23576 33876 23588
rect 33735 23548 33876 23576
rect 33735 23545 33747 23548
rect 33689 23539 33747 23545
rect 33870 23536 33876 23548
rect 33928 23536 33934 23588
rect 27856 23480 28488 23508
rect 28905 23511 28963 23517
rect 27856 23468 27862 23480
rect 28905 23477 28917 23511
rect 28951 23508 28963 23511
rect 31110 23508 31116 23520
rect 28951 23480 31116 23508
rect 28951 23477 28963 23480
rect 28905 23471 28963 23477
rect 31110 23468 31116 23480
rect 31168 23468 31174 23520
rect 31386 23468 31392 23520
rect 31444 23468 31450 23520
rect 31846 23468 31852 23520
rect 31904 23468 31910 23520
rect 32214 23468 32220 23520
rect 32272 23508 32278 23520
rect 33229 23511 33287 23517
rect 33229 23508 33241 23511
rect 32272 23480 33241 23508
rect 32272 23468 32278 23480
rect 33229 23477 33241 23480
rect 33275 23477 33287 23511
rect 33229 23471 33287 23477
rect 33778 23468 33784 23520
rect 33836 23468 33842 23520
rect 34348 23508 34376 23604
rect 35618 23536 35624 23588
rect 35676 23576 35682 23588
rect 38105 23579 38163 23585
rect 38105 23576 38117 23579
rect 35676 23548 38117 23576
rect 35676 23536 35682 23548
rect 38105 23545 38117 23548
rect 38151 23545 38163 23579
rect 38105 23539 38163 23545
rect 38286 23536 38292 23588
rect 38344 23576 38350 23588
rect 41785 23579 41843 23585
rect 41785 23576 41797 23579
rect 38344 23548 41797 23576
rect 38344 23536 38350 23548
rect 41785 23545 41797 23548
rect 41831 23545 41843 23579
rect 41785 23539 41843 23545
rect 43438 23536 43444 23588
rect 43496 23576 43502 23588
rect 44453 23579 44511 23585
rect 44453 23576 44465 23579
rect 43496 23548 44465 23576
rect 43496 23536 43502 23548
rect 44453 23545 44465 23548
rect 44499 23545 44511 23579
rect 44453 23539 44511 23545
rect 39301 23511 39359 23517
rect 39301 23508 39313 23511
rect 34348 23480 39313 23508
rect 39301 23477 39313 23480
rect 39347 23477 39359 23511
rect 39301 23471 39359 23477
rect 40218 23468 40224 23520
rect 40276 23508 40282 23520
rect 41046 23508 41052 23520
rect 40276 23480 41052 23508
rect 40276 23468 40282 23480
rect 41046 23468 41052 23480
rect 41104 23468 41110 23520
rect 43714 23468 43720 23520
rect 43772 23468 43778 23520
rect 46934 23468 46940 23520
rect 46992 23468 46998 23520
rect 48682 23468 48688 23520
rect 48740 23468 48746 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 2746 23276 14473 23304
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 2746 23100 2774 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 16206 23264 16212 23316
rect 16264 23304 16270 23316
rect 18966 23304 18972 23316
rect 16264 23276 18972 23304
rect 16264 23264 16270 23276
rect 18966 23264 18972 23276
rect 19024 23264 19030 23316
rect 23014 23304 23020 23316
rect 19306 23276 23020 23304
rect 3421 23239 3479 23245
rect 3421 23205 3433 23239
rect 3467 23236 3479 23239
rect 6822 23236 6828 23248
rect 3467 23208 6828 23236
rect 3467 23205 3479 23208
rect 3421 23199 3479 23205
rect 6822 23196 6828 23208
rect 6880 23196 6886 23248
rect 9122 23196 9128 23248
rect 9180 23196 9186 23248
rect 11146 23196 11152 23248
rect 11204 23196 11210 23248
rect 18877 23239 18935 23245
rect 18877 23205 18889 23239
rect 18923 23236 18935 23239
rect 19306 23236 19334 23276
rect 23014 23264 23020 23276
rect 23072 23264 23078 23316
rect 23106 23264 23112 23316
rect 23164 23304 23170 23316
rect 25777 23307 25835 23313
rect 25777 23304 25789 23307
rect 23164 23276 25789 23304
rect 23164 23264 23170 23276
rect 25777 23273 25789 23276
rect 25823 23273 25835 23307
rect 28997 23307 29055 23313
rect 28997 23304 29009 23307
rect 25777 23267 25835 23273
rect 26160 23276 29009 23304
rect 18923 23208 19334 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 21818 23196 21824 23248
rect 21876 23196 21882 23248
rect 24670 23196 24676 23248
rect 24728 23196 24734 23248
rect 3605 23171 3663 23177
rect 3605 23137 3617 23171
rect 3651 23168 3663 23171
rect 5534 23168 5540 23180
rect 3651 23140 5540 23168
rect 3651 23137 3663 23140
rect 3605 23131 3663 23137
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11164 23168 11192 23196
rect 7944 23140 11192 23168
rect 11701 23171 11759 23177
rect 1811 23072 2774 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 3970 23060 3976 23112
rect 4028 23060 4034 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 5368 23032 5396 23063
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 7064 23072 7205 23100
rect 7064 23060 7070 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 7374 23060 7380 23112
rect 7432 23100 7438 23112
rect 7944 23100 7972 23140
rect 11701 23137 11713 23171
rect 11747 23168 11759 23171
rect 12526 23168 12532 23180
rect 11747 23140 12532 23168
rect 11747 23137 11759 23140
rect 11701 23131 11759 23137
rect 12526 23128 12532 23140
rect 12584 23128 12590 23180
rect 17954 23168 17960 23180
rect 15488 23140 17960 23168
rect 7432 23072 7972 23100
rect 7432 23060 7438 23072
rect 9398 23060 9404 23112
rect 9456 23060 9462 23112
rect 14369 23103 14427 23109
rect 14369 23069 14381 23103
rect 14415 23100 14427 23103
rect 14550 23100 14556 23112
rect 14415 23072 14556 23100
rect 14415 23069 14427 23072
rect 14369 23063 14427 23069
rect 14550 23060 14556 23072
rect 14608 23060 14614 23112
rect 15488 23109 15516 23140
rect 17954 23128 17960 23140
rect 18012 23128 18018 23180
rect 19702 23128 19708 23180
rect 19760 23168 19766 23180
rect 20073 23171 20131 23177
rect 20073 23168 20085 23171
rect 19760 23140 20085 23168
rect 19760 23128 19766 23140
rect 20073 23137 20085 23140
rect 20119 23168 20131 23171
rect 20346 23168 20352 23180
rect 20119 23140 20352 23168
rect 20119 23137 20131 23140
rect 20073 23131 20131 23137
rect 20346 23128 20352 23140
rect 20404 23128 20410 23180
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 20496 23140 21496 23168
rect 20496 23128 20502 23140
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 21468 23086 21496 23140
rect 22278 23128 22284 23180
rect 22336 23168 22342 23180
rect 23290 23168 23296 23180
rect 22336 23140 23296 23168
rect 22336 23128 22342 23140
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23566 23128 23572 23180
rect 23624 23168 23630 23180
rect 23750 23168 23756 23180
rect 23624 23140 23756 23168
rect 23624 23128 23630 23140
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 26160 23168 26188 23276
rect 28997 23273 29009 23276
rect 29043 23304 29055 23307
rect 30098 23304 30104 23316
rect 29043 23276 30104 23304
rect 29043 23273 29055 23276
rect 28997 23267 29055 23273
rect 30098 23264 30104 23276
rect 30156 23264 30162 23316
rect 30190 23264 30196 23316
rect 30248 23304 30254 23316
rect 30248 23276 32628 23304
rect 30248 23264 30254 23276
rect 28534 23196 28540 23248
rect 28592 23236 28598 23248
rect 29086 23236 29092 23248
rect 28592 23208 29092 23236
rect 28592 23196 28598 23208
rect 29086 23196 29092 23208
rect 29144 23196 29150 23248
rect 32600 23236 32628 23276
rect 32766 23264 32772 23316
rect 32824 23304 32830 23316
rect 34885 23307 34943 23313
rect 34885 23304 34897 23307
rect 32824 23276 34897 23304
rect 32824 23264 32830 23276
rect 34885 23273 34897 23276
rect 34931 23273 34943 23307
rect 34885 23267 34943 23273
rect 34974 23264 34980 23316
rect 35032 23304 35038 23316
rect 36998 23304 37004 23316
rect 35032 23276 37004 23304
rect 35032 23264 35038 23276
rect 36998 23264 37004 23276
rect 37056 23264 37062 23316
rect 37090 23264 37096 23316
rect 37148 23304 37154 23316
rect 37148 23276 40816 23304
rect 37148 23264 37154 23276
rect 34149 23239 34207 23245
rect 34149 23236 34161 23239
rect 32600 23208 34161 23236
rect 34149 23205 34161 23208
rect 34195 23205 34207 23239
rect 34149 23199 34207 23205
rect 34238 23196 34244 23248
rect 34296 23236 34302 23248
rect 36446 23236 36452 23248
rect 34296 23208 36452 23236
rect 34296 23196 34302 23208
rect 36446 23196 36452 23208
rect 36504 23236 36510 23248
rect 36817 23239 36875 23245
rect 36504 23208 36676 23236
rect 36504 23196 36510 23208
rect 25271 23140 26188 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 26418 23128 26424 23180
rect 26476 23128 26482 23180
rect 27246 23128 27252 23180
rect 27304 23168 27310 23180
rect 28902 23168 28908 23180
rect 27304 23140 28908 23168
rect 27304 23128 27310 23140
rect 28902 23128 28908 23140
rect 28960 23168 28966 23180
rect 29273 23171 29331 23177
rect 29273 23168 29285 23171
rect 28960 23140 29285 23168
rect 28960 23128 28966 23140
rect 29273 23137 29285 23140
rect 29319 23168 29331 23171
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 29319 23140 29745 23168
rect 29319 23137 29331 23140
rect 29273 23131 29331 23137
rect 29733 23137 29745 23140
rect 29779 23137 29791 23171
rect 29733 23131 29791 23137
rect 30006 23128 30012 23180
rect 30064 23128 30070 23180
rect 32582 23128 32588 23180
rect 32640 23168 32646 23180
rect 32640 23140 34376 23168
rect 32640 23128 32646 23140
rect 34348 23112 34376 23140
rect 34790 23128 34796 23180
rect 34848 23168 34854 23180
rect 34848 23140 35664 23168
rect 34848 23128 34854 23140
rect 23842 23060 23848 23112
rect 23900 23100 23906 23112
rect 26050 23100 26056 23112
rect 23900 23072 26056 23100
rect 23900 23060 23906 23072
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 26200 23072 26249 23100
rect 26200 23060 26206 23072
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 31754 23100 31760 23112
rect 31142 23072 31760 23100
rect 26237 23063 26295 23069
rect 31754 23060 31760 23072
rect 31812 23060 31818 23112
rect 31938 23060 31944 23112
rect 31996 23060 32002 23112
rect 32030 23060 32036 23112
rect 32088 23100 32094 23112
rect 32950 23100 32956 23112
rect 32088 23072 32956 23100
rect 32088 23060 32094 23072
rect 32950 23060 32956 23072
rect 33008 23060 33014 23112
rect 33045 23103 33103 23109
rect 33045 23069 33057 23103
rect 33091 23069 33103 23103
rect 33045 23063 33103 23069
rect 3252 23004 5396 23032
rect 934 22924 940 22976
rect 992 22964 998 22976
rect 3252 22964 3280 23004
rect 5626 22992 5632 23044
rect 5684 23032 5690 23044
rect 5684 23004 6592 23032
rect 5684 22992 5690 23004
rect 992 22936 3280 22964
rect 4203 22967 4261 22973
rect 992 22924 998 22936
rect 4203 22933 4215 22967
rect 4249 22964 4261 22967
rect 6454 22964 6460 22976
rect 4249 22936 6460 22964
rect 4249 22933 4261 22936
rect 4203 22927 4261 22933
rect 6454 22924 6460 22936
rect 6512 22924 6518 22976
rect 6564 22964 6592 23004
rect 9674 22992 9680 23044
rect 9732 22992 9738 23044
rect 11422 23032 11428 23044
rect 10902 23004 11428 23032
rect 11422 22992 11428 23004
rect 11480 23032 11486 23044
rect 11698 23032 11704 23044
rect 11480 23004 11704 23032
rect 11480 22992 11486 23004
rect 11698 22992 11704 23004
rect 11756 22992 11762 23044
rect 11977 23035 12035 23041
rect 11977 23001 11989 23035
rect 12023 23032 12035 23035
rect 12066 23032 12072 23044
rect 12023 23004 12072 23032
rect 12023 23001 12035 23004
rect 11977 22995 12035 23001
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 13814 23032 13820 23044
rect 13202 23004 13820 23032
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 16485 23035 16543 23041
rect 16485 23001 16497 23035
rect 16531 23032 16543 23035
rect 17310 23032 17316 23044
rect 16531 23004 17316 23032
rect 16531 23001 16543 23004
rect 16485 22995 16543 23001
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 17402 22992 17408 23044
rect 17460 22992 17466 23044
rect 18414 22992 18420 23044
rect 18472 22992 18478 23044
rect 20349 23035 20407 23041
rect 20349 23001 20361 23035
rect 20395 23032 20407 23035
rect 20622 23032 20628 23044
rect 20395 23004 20628 23032
rect 20395 23001 20407 23004
rect 20349 22995 20407 23001
rect 20622 22992 20628 23004
rect 20680 22992 20686 23044
rect 21652 23004 22094 23032
rect 12618 22964 12624 22976
rect 6564 22936 12624 22964
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 13449 22967 13507 22973
rect 13449 22964 13461 22967
rect 12768 22936 13461 22964
rect 12768 22924 12774 22936
rect 13449 22933 13461 22936
rect 13495 22933 13507 22967
rect 13449 22927 13507 22933
rect 14550 22924 14556 22976
rect 14608 22964 14614 22976
rect 14921 22967 14979 22973
rect 14921 22964 14933 22967
rect 14608 22936 14933 22964
rect 14608 22924 14614 22936
rect 14921 22933 14933 22936
rect 14967 22933 14979 22967
rect 14921 22927 14979 22933
rect 16298 22924 16304 22976
rect 16356 22964 16362 22976
rect 18322 22964 18328 22976
rect 16356 22936 18328 22964
rect 16356 22924 16362 22936
rect 18322 22924 18328 22936
rect 18380 22924 18386 22976
rect 19429 22967 19487 22973
rect 19429 22933 19441 22967
rect 19475 22964 19487 22967
rect 21652 22964 21680 23004
rect 19475 22936 21680 22964
rect 22066 22964 22094 23004
rect 22554 22992 22560 23044
rect 22612 22992 22618 23044
rect 23566 22992 23572 23044
rect 23624 22992 23630 23044
rect 24949 23035 25007 23041
rect 24949 23032 24961 23035
rect 23860 23004 24961 23032
rect 23860 22964 23888 23004
rect 24949 23001 24961 23004
rect 24995 23001 25007 23035
rect 24949 22995 25007 23001
rect 26326 22992 26332 23044
rect 26384 23032 26390 23044
rect 26789 23035 26847 23041
rect 26789 23032 26801 23035
rect 26384 23004 26801 23032
rect 26384 22992 26390 23004
rect 26789 23001 26801 23004
rect 26835 23001 26847 23035
rect 26789 22995 26847 23001
rect 27430 22992 27436 23044
rect 27488 23032 27494 23044
rect 27525 23035 27583 23041
rect 27525 23032 27537 23035
rect 27488 23004 27537 23032
rect 27488 22992 27494 23004
rect 27525 23001 27537 23004
rect 27571 23001 27583 23035
rect 29086 23032 29092 23044
rect 28750 23004 29092 23032
rect 27525 22995 27583 23001
rect 29086 22992 29092 23004
rect 29144 22992 29150 23044
rect 33060 23032 33088 23063
rect 34330 23060 34336 23112
rect 34388 23060 34394 23112
rect 35066 23060 35072 23112
rect 35124 23060 35130 23112
rect 35526 23060 35532 23112
rect 35584 23060 35590 23112
rect 35636 23100 35664 23140
rect 35710 23128 35716 23180
rect 35768 23168 35774 23180
rect 36648 23168 36676 23208
rect 36817 23205 36829 23239
rect 36863 23236 36875 23239
rect 36906 23236 36912 23248
rect 36863 23208 36912 23236
rect 36863 23205 36875 23208
rect 36817 23199 36875 23205
rect 36906 23196 36912 23208
rect 36964 23196 36970 23248
rect 37274 23196 37280 23248
rect 37332 23236 37338 23248
rect 40681 23239 40739 23245
rect 40681 23236 40693 23239
rect 37332 23208 40693 23236
rect 37332 23196 37338 23208
rect 40681 23205 40693 23208
rect 40727 23205 40739 23239
rect 40681 23199 40739 23205
rect 36722 23168 36728 23180
rect 35768 23140 36584 23168
rect 36648 23140 36728 23168
rect 35768 23128 35774 23140
rect 35805 23103 35863 23109
rect 35805 23100 35817 23103
rect 35636 23072 35817 23100
rect 35805 23069 35817 23072
rect 35851 23069 35863 23103
rect 36556 23100 36584 23140
rect 36722 23128 36728 23140
rect 36780 23128 36786 23180
rect 39485 23171 39543 23177
rect 39485 23168 39497 23171
rect 36832 23140 39497 23168
rect 36832 23100 36860 23140
rect 39485 23137 39497 23140
rect 39531 23137 39543 23171
rect 40788 23168 40816 23276
rect 40862 23196 40868 23248
rect 40920 23236 40926 23248
rect 40920 23208 41414 23236
rect 40920 23196 40926 23208
rect 41386 23168 41414 23208
rect 42429 23171 42487 23177
rect 42429 23168 42441 23171
rect 40788 23140 41000 23168
rect 41386 23140 42441 23168
rect 39485 23131 39543 23137
rect 36556 23072 36860 23100
rect 35805 23063 35863 23069
rect 36998 23060 37004 23112
rect 37056 23100 37062 23112
rect 37458 23100 37464 23112
rect 37056 23072 37464 23100
rect 37056 23060 37062 23072
rect 37458 23060 37464 23072
rect 37516 23060 37522 23112
rect 38470 23060 38476 23112
rect 38528 23060 38534 23112
rect 38930 23060 38936 23112
rect 38988 23060 38994 23112
rect 39758 23060 39764 23112
rect 39816 23100 39822 23112
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 39816 23072 40233 23100
rect 39816 23060 39822 23072
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 40221 23063 40279 23069
rect 40862 23060 40868 23112
rect 40920 23060 40926 23112
rect 40972 23100 41000 23140
rect 41138 23100 41144 23112
rect 40972 23072 41144 23100
rect 41138 23060 41144 23072
rect 41196 23100 41202 23112
rect 42168 23109 42196 23140
rect 42429 23137 42441 23140
rect 42475 23137 42487 23171
rect 42429 23131 42487 23137
rect 41509 23103 41567 23109
rect 41509 23100 41521 23103
rect 41196 23072 41521 23100
rect 41196 23060 41202 23072
rect 41509 23069 41521 23072
rect 41555 23069 41567 23103
rect 41509 23063 41567 23069
rect 42153 23103 42211 23109
rect 42153 23069 42165 23103
rect 42199 23069 42211 23103
rect 42153 23063 42211 23069
rect 34974 23032 34980 23044
rect 31496 23004 33088 23032
rect 33612 23004 34980 23032
rect 22066 22936 23888 22964
rect 19475 22933 19487 22936
rect 19429 22927 19487 22933
rect 24026 22924 24032 22976
rect 24084 22924 24090 22976
rect 25130 22924 25136 22976
rect 25188 22924 25194 22976
rect 25682 22924 25688 22976
rect 25740 22964 25746 22976
rect 25958 22964 25964 22976
rect 25740 22936 25964 22964
rect 25740 22924 25746 22936
rect 25958 22924 25964 22936
rect 26016 22964 26022 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 26016 22936 26157 22964
rect 26016 22924 26022 22936
rect 26145 22933 26157 22936
rect 26191 22964 26203 22967
rect 26418 22964 26424 22976
rect 26191 22936 26424 22964
rect 26191 22933 26203 22936
rect 26145 22927 26203 22933
rect 26418 22924 26424 22936
rect 26476 22924 26482 22976
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 30374 22964 30380 22976
rect 27764 22936 30380 22964
rect 27764 22924 27770 22936
rect 30374 22924 30380 22936
rect 30432 22924 30438 22976
rect 30650 22924 30656 22976
rect 30708 22964 30714 22976
rect 31496 22973 31524 23004
rect 31481 22967 31539 22973
rect 31481 22964 31493 22967
rect 30708 22936 31493 22964
rect 30708 22924 30714 22936
rect 31481 22933 31493 22936
rect 31527 22933 31539 22967
rect 31481 22927 31539 22933
rect 31570 22924 31576 22976
rect 31628 22964 31634 22976
rect 32585 22967 32643 22973
rect 32585 22964 32597 22967
rect 31628 22936 32597 22964
rect 31628 22924 31634 22936
rect 32585 22933 32597 22936
rect 32631 22933 32643 22967
rect 32585 22927 32643 22933
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 33612 22964 33640 23004
rect 34974 22992 34980 23004
rect 35032 22992 35038 23044
rect 35158 22992 35164 23044
rect 35216 23032 35222 23044
rect 37366 23032 37372 23044
rect 35216 23004 37372 23032
rect 35216 22992 35222 23004
rect 37366 22992 37372 23004
rect 37424 22992 37430 23044
rect 37550 22992 37556 23044
rect 37608 22992 37614 23044
rect 38286 22992 38292 23044
rect 38344 22992 38350 23044
rect 39574 22992 39580 23044
rect 39632 23032 39638 23044
rect 39632 23004 41368 23032
rect 39632 22992 39638 23004
rect 33008 22936 33640 22964
rect 33008 22924 33014 22936
rect 33686 22924 33692 22976
rect 33744 22924 33750 22976
rect 35894 22924 35900 22976
rect 35952 22964 35958 22976
rect 37182 22964 37188 22976
rect 35952 22936 37188 22964
rect 35952 22924 35958 22936
rect 37182 22924 37188 22936
rect 37240 22924 37246 22976
rect 37642 22924 37648 22976
rect 37700 22924 37706 22976
rect 39114 22924 39120 22976
rect 39172 22924 39178 22976
rect 39850 22924 39856 22976
rect 39908 22964 39914 22976
rect 41340 22973 41368 23004
rect 40037 22967 40095 22973
rect 40037 22964 40049 22967
rect 39908 22936 40049 22964
rect 39908 22924 39914 22936
rect 40037 22933 40049 22936
rect 40083 22933 40095 22967
rect 40037 22927 40095 22933
rect 41325 22967 41383 22973
rect 41325 22933 41337 22967
rect 41371 22933 41383 22967
rect 41325 22927 41383 22933
rect 41966 22924 41972 22976
rect 42024 22924 42030 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 658 22720 664 22772
rect 716 22760 722 22772
rect 716 22732 7972 22760
rect 716 22720 722 22732
rect 5166 22692 5172 22704
rect 3528 22664 5172 22692
rect 3528 22633 3556 22664
rect 5166 22652 5172 22664
rect 5224 22652 5230 22704
rect 5258 22652 5264 22704
rect 5316 22692 5322 22704
rect 5537 22695 5595 22701
rect 5537 22692 5549 22695
rect 5316 22664 5549 22692
rect 5316 22652 5322 22664
rect 5537 22661 5549 22664
rect 5583 22661 5595 22695
rect 5537 22655 5595 22661
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22692 6699 22695
rect 7098 22692 7104 22704
rect 6687 22664 7104 22692
rect 6687 22661 6699 22664
rect 6641 22655 6699 22661
rect 7098 22652 7104 22664
rect 7156 22652 7162 22704
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 3513 22627 3571 22633
rect 1811 22596 3464 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3436 22420 3464 22596
rect 3513 22593 3525 22627
rect 3559 22593 3571 22627
rect 3513 22587 3571 22593
rect 4614 22584 4620 22636
rect 4672 22584 4678 22636
rect 6914 22624 6920 22636
rect 5000 22596 6920 22624
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 5000 22556 5028 22596
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7944 22633 7972 22732
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 11054 22760 11060 22772
rect 9732 22732 11060 22760
rect 9732 22720 9738 22732
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 12526 22720 12532 22772
rect 12584 22720 12590 22772
rect 12618 22720 12624 22772
rect 12676 22760 12682 22772
rect 14826 22760 14832 22772
rect 12676 22732 14832 22760
rect 12676 22720 12682 22732
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 18601 22763 18659 22769
rect 15028 22732 18552 22760
rect 8570 22652 8576 22704
rect 8628 22692 8634 22704
rect 8628 22664 9904 22692
rect 8628 22652 8634 22664
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22624 7251 22627
rect 7929 22627 7987 22633
rect 7239 22596 7880 22624
rect 7239 22593 7251 22596
rect 7193 22587 7251 22593
rect 4203 22528 5028 22556
rect 5184 22528 6868 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 5184 22420 5212 22528
rect 5258 22448 5264 22500
rect 5316 22488 5322 22500
rect 6733 22491 6791 22497
rect 6733 22488 6745 22491
rect 5316 22460 6745 22488
rect 5316 22448 5322 22460
rect 6733 22457 6745 22460
rect 6779 22457 6791 22491
rect 6840 22488 6868 22528
rect 7374 22516 7380 22568
rect 7432 22516 7438 22568
rect 7852 22556 7880 22596
rect 7929 22593 7941 22627
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 8588 22596 9720 22624
rect 8588 22556 8616 22596
rect 7852 22528 8616 22556
rect 8662 22516 8668 22568
rect 8720 22516 8726 22568
rect 9692 22556 9720 22596
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 9876 22624 9904 22664
rect 10686 22652 10692 22704
rect 10744 22652 10750 22704
rect 11790 22652 11796 22704
rect 11848 22652 11854 22704
rect 12544 22692 12572 22720
rect 12452 22664 12572 22692
rect 11330 22624 11336 22636
rect 9876 22596 11336 22624
rect 11330 22584 11336 22596
rect 11388 22584 11394 22636
rect 12452 22633 12480 22664
rect 12710 22652 12716 22704
rect 12768 22652 12774 22704
rect 12437 22627 12495 22633
rect 12437 22593 12449 22627
rect 12483 22593 12495 22627
rect 12437 22587 12495 22593
rect 13814 22584 13820 22636
rect 13872 22584 13878 22636
rect 14918 22584 14924 22636
rect 14976 22584 14982 22636
rect 10962 22556 10968 22568
rect 9692 22528 10968 22556
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 11146 22516 11152 22568
rect 11204 22556 11210 22568
rect 15028 22556 15056 22732
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 16761 22695 16819 22701
rect 16761 22661 16773 22695
rect 16807 22692 16819 22695
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16807 22664 17141 22692
rect 16807 22661 16819 22664
rect 16761 22655 16819 22661
rect 17129 22661 17141 22664
rect 17175 22692 17187 22695
rect 17218 22692 17224 22704
rect 17175 22664 17224 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 18414 22692 18420 22704
rect 18354 22664 18420 22692
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 18524 22692 18552 22732
rect 18601 22729 18613 22763
rect 18647 22760 18659 22763
rect 18874 22760 18880 22772
rect 18647 22732 18880 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 19061 22763 19119 22769
rect 19061 22729 19073 22763
rect 19107 22760 19119 22763
rect 24857 22763 24915 22769
rect 24857 22760 24869 22763
rect 19107 22732 21312 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19518 22692 19524 22704
rect 18524 22664 19524 22692
rect 19518 22652 19524 22664
rect 19576 22652 19582 22704
rect 19978 22652 19984 22704
rect 20036 22652 20042 22704
rect 20438 22652 20444 22704
rect 20496 22652 20502 22704
rect 19702 22584 19708 22636
rect 19760 22584 19766 22636
rect 11204 22528 15056 22556
rect 16853 22559 16911 22565
rect 11204 22516 11210 22528
rect 16853 22525 16865 22559
rect 16899 22525 16911 22559
rect 21284 22556 21312 22732
rect 22020 22732 24869 22760
rect 22020 22633 22048 22732
rect 24857 22729 24869 22732
rect 24903 22729 24915 22763
rect 24857 22723 24915 22729
rect 25685 22763 25743 22769
rect 25685 22729 25697 22763
rect 25731 22760 25743 22763
rect 26326 22760 26332 22772
rect 25731 22732 26332 22760
rect 25731 22729 25743 22732
rect 25685 22723 25743 22729
rect 23290 22692 23296 22704
rect 23124 22664 23296 22692
rect 23124 22633 23152 22664
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 23385 22695 23443 22701
rect 23385 22661 23397 22695
rect 23431 22692 23443 22695
rect 23474 22692 23480 22704
rect 23431 22664 23480 22692
rect 23431 22661 23443 22664
rect 23385 22655 23443 22661
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 23842 22652 23848 22704
rect 23900 22652 23906 22704
rect 24872 22692 24900 22723
rect 26326 22720 26332 22732
rect 26384 22720 26390 22772
rect 26789 22763 26847 22769
rect 26789 22729 26801 22763
rect 26835 22760 26847 22763
rect 27246 22760 27252 22772
rect 26835 22732 27252 22760
rect 26835 22729 26847 22732
rect 26789 22723 26847 22729
rect 27246 22720 27252 22732
rect 27304 22720 27310 22772
rect 28902 22720 28908 22772
rect 28960 22760 28966 22772
rect 31570 22760 31576 22772
rect 28960 22732 31576 22760
rect 28960 22720 28966 22732
rect 31570 22720 31576 22732
rect 31628 22720 31634 22772
rect 31662 22720 31668 22772
rect 31720 22760 31726 22772
rect 32953 22763 33011 22769
rect 32953 22760 32965 22763
rect 31720 22732 32965 22760
rect 31720 22720 31726 22732
rect 32953 22729 32965 22732
rect 32999 22729 33011 22763
rect 32953 22723 33011 22729
rect 33226 22720 33232 22772
rect 33284 22760 33290 22772
rect 33321 22763 33379 22769
rect 33321 22760 33333 22763
rect 33284 22732 33333 22760
rect 33284 22720 33290 22732
rect 33321 22729 33333 22732
rect 33367 22760 33379 22763
rect 33870 22760 33876 22772
rect 33367 22732 33876 22760
rect 33367 22729 33379 22732
rect 33321 22723 33379 22729
rect 33870 22720 33876 22732
rect 33928 22760 33934 22772
rect 33928 22732 34284 22760
rect 33928 22720 33934 22732
rect 24872 22664 25912 22692
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 22738 22556 22744 22568
rect 21284 22528 22744 22556
rect 16853 22519 16911 22525
rect 11977 22491 12035 22497
rect 11977 22488 11989 22491
rect 6840 22460 11989 22488
rect 6733 22451 6791 22457
rect 11977 22457 11989 22460
rect 12023 22457 12035 22491
rect 16758 22488 16764 22500
rect 11977 22451 12035 22457
rect 14108 22460 16764 22488
rect 3436 22392 5212 22420
rect 5534 22380 5540 22432
rect 5592 22420 5598 22432
rect 6454 22420 6460 22432
rect 5592 22392 6460 22420
rect 5592 22380 5598 22392
rect 6454 22380 6460 22392
rect 6512 22380 6518 22432
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 14108 22420 14136 22460
rect 16758 22448 16764 22460
rect 16816 22448 16822 22500
rect 11112 22392 14136 22420
rect 11112 22380 11118 22392
rect 14182 22380 14188 22432
rect 14240 22380 14246 22432
rect 14550 22380 14556 22432
rect 14608 22380 14614 22432
rect 16868 22420 16896 22519
rect 22738 22516 22744 22528
rect 22796 22516 22802 22568
rect 23014 22516 23020 22568
rect 23072 22556 23078 22568
rect 25222 22556 25228 22568
rect 23072 22528 25228 22556
rect 23072 22516 23078 22528
rect 25222 22516 25228 22528
rect 25280 22516 25286 22568
rect 25884 22565 25912 22664
rect 27157 22627 27215 22633
rect 27157 22593 27169 22627
rect 27203 22593 27215 22627
rect 27264 22624 27292 22720
rect 30098 22692 30104 22704
rect 29854 22664 30104 22692
rect 30098 22652 30104 22664
rect 30156 22652 30162 22704
rect 33686 22692 33692 22704
rect 30208 22664 33692 22692
rect 28353 22627 28411 22633
rect 28353 22624 28365 22627
rect 27264 22596 28365 22624
rect 27157 22587 27215 22593
rect 28353 22593 28365 22596
rect 28399 22593 28411 22627
rect 28353 22587 28411 22593
rect 25777 22559 25835 22565
rect 25777 22525 25789 22559
rect 25823 22525 25835 22559
rect 25777 22519 25835 22525
rect 25869 22559 25927 22565
rect 25869 22525 25881 22559
rect 25915 22525 25927 22559
rect 27172 22556 27200 22587
rect 27246 22556 27252 22568
rect 25869 22519 25927 22525
rect 25976 22528 27108 22556
rect 27172 22528 27252 22556
rect 23106 22488 23112 22500
rect 21008 22460 23112 22488
rect 17126 22420 17132 22432
rect 16868 22392 17132 22420
rect 17126 22380 17132 22392
rect 17184 22420 17190 22432
rect 18506 22420 18512 22432
rect 17184 22392 18512 22420
rect 17184 22380 17190 22392
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 18966 22380 18972 22432
rect 19024 22420 19030 22432
rect 21008 22420 21036 22460
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 25682 22488 25688 22500
rect 25240 22460 25688 22488
rect 19024 22392 21036 22420
rect 19024 22380 19030 22392
rect 21450 22380 21456 22432
rect 21508 22380 21514 22432
rect 22649 22423 22707 22429
rect 22649 22389 22661 22423
rect 22695 22420 22707 22423
rect 23566 22420 23572 22432
rect 22695 22392 23572 22420
rect 22695 22389 22707 22392
rect 22649 22383 22707 22389
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 23750 22380 23756 22432
rect 23808 22420 23814 22432
rect 25240 22420 25268 22460
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 25792 22488 25820 22519
rect 25976 22488 26004 22528
rect 25792 22460 26004 22488
rect 26050 22448 26056 22500
rect 26108 22488 26114 22500
rect 26329 22491 26387 22497
rect 26329 22488 26341 22491
rect 26108 22460 26341 22488
rect 26108 22448 26114 22460
rect 26329 22457 26341 22460
rect 26375 22457 26387 22491
rect 27080 22488 27108 22528
rect 27246 22516 27252 22528
rect 27304 22516 27310 22568
rect 28629 22559 28687 22565
rect 28629 22525 28641 22559
rect 28675 22556 28687 22559
rect 30208 22556 30236 22664
rect 33686 22652 33692 22664
rect 33744 22652 33750 22704
rect 34256 22692 34284 22732
rect 34330 22720 34336 22772
rect 34388 22760 34394 22772
rect 37461 22763 37519 22769
rect 37461 22760 37473 22763
rect 34388 22732 37473 22760
rect 34388 22720 34394 22732
rect 37461 22729 37473 22732
rect 37507 22729 37519 22763
rect 39945 22763 40003 22769
rect 39945 22760 39957 22763
rect 37461 22723 37519 22729
rect 37568 22732 39957 22760
rect 34422 22692 34428 22704
rect 34256 22664 34428 22692
rect 34422 22652 34428 22664
rect 34480 22652 34486 22704
rect 36630 22652 36636 22704
rect 36688 22692 36694 22704
rect 37277 22695 37335 22701
rect 37277 22692 37289 22695
rect 36688 22664 37289 22692
rect 36688 22652 36694 22664
rect 37277 22661 37289 22664
rect 37323 22661 37335 22695
rect 37277 22655 37335 22661
rect 37366 22652 37372 22704
rect 37424 22692 37430 22704
rect 37568 22692 37596 22732
rect 39945 22729 39957 22732
rect 39991 22729 40003 22763
rect 39945 22723 40003 22729
rect 40034 22720 40040 22772
rect 40092 22760 40098 22772
rect 40129 22763 40187 22769
rect 40129 22760 40141 22763
rect 40092 22732 40141 22760
rect 40092 22720 40098 22732
rect 40129 22729 40141 22732
rect 40175 22729 40187 22763
rect 40129 22723 40187 22729
rect 41138 22720 41144 22772
rect 41196 22720 41202 22772
rect 39482 22692 39488 22704
rect 37424 22664 37596 22692
rect 39422 22664 39488 22692
rect 37424 22652 37430 22664
rect 39482 22652 39488 22664
rect 39540 22692 39546 22704
rect 40405 22695 40463 22701
rect 40405 22692 40417 22695
rect 39540 22664 40417 22692
rect 39540 22652 39546 22664
rect 40405 22661 40417 22664
rect 40451 22692 40463 22695
rect 43898 22692 43904 22704
rect 40451 22664 43904 22692
rect 40451 22661 40463 22664
rect 40405 22655 40463 22661
rect 43898 22652 43904 22664
rect 43956 22652 43962 22704
rect 30929 22627 30987 22633
rect 30929 22593 30941 22627
rect 30975 22624 30987 22627
rect 31202 22624 31208 22636
rect 30975 22596 31208 22624
rect 30975 22593 30987 22596
rect 30929 22587 30987 22593
rect 31202 22584 31208 22596
rect 31260 22584 31266 22636
rect 31846 22584 31852 22636
rect 31904 22584 31910 22636
rect 32306 22584 32312 22636
rect 32364 22584 32370 22636
rect 33870 22584 33876 22636
rect 33928 22584 33934 22636
rect 34609 22627 34667 22633
rect 34609 22593 34621 22627
rect 34655 22624 34667 22627
rect 34698 22624 34704 22636
rect 34655 22596 34704 22624
rect 34655 22593 34667 22596
rect 34609 22587 34667 22593
rect 34698 22584 34704 22596
rect 34756 22584 34762 22636
rect 35618 22584 35624 22636
rect 35676 22624 35682 22636
rect 35713 22627 35771 22633
rect 35713 22624 35725 22627
rect 35676 22596 35725 22624
rect 35676 22584 35682 22596
rect 35713 22593 35725 22596
rect 35759 22593 35771 22627
rect 35713 22587 35771 22593
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22624 36507 22627
rect 36722 22624 36728 22636
rect 36495 22596 36728 22624
rect 36495 22593 36507 22596
rect 36449 22587 36507 22593
rect 36722 22584 36728 22596
rect 36780 22584 36786 22636
rect 36832 22596 37964 22624
rect 28675 22528 30236 22556
rect 28675 22525 28687 22528
rect 28629 22519 28687 22525
rect 31018 22516 31024 22568
rect 31076 22516 31082 22568
rect 31110 22516 31116 22568
rect 31168 22516 31174 22568
rect 31570 22516 31576 22568
rect 31628 22556 31634 22568
rect 33778 22556 33784 22568
rect 31628 22528 33784 22556
rect 31628 22516 31634 22528
rect 33778 22516 33784 22528
rect 33836 22516 33842 22568
rect 34330 22516 34336 22568
rect 34388 22516 34394 22568
rect 35897 22559 35955 22565
rect 35897 22525 35909 22559
rect 35943 22556 35955 22559
rect 35986 22556 35992 22568
rect 35943 22528 35992 22556
rect 35943 22525 35955 22528
rect 35897 22519 35955 22525
rect 35986 22516 35992 22528
rect 36044 22516 36050 22568
rect 27614 22488 27620 22500
rect 27080 22460 27620 22488
rect 26329 22451 26387 22457
rect 27614 22448 27620 22460
rect 27672 22448 27678 22500
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 30561 22491 30619 22497
rect 30561 22488 30573 22491
rect 30432 22460 30573 22488
rect 30432 22448 30438 22460
rect 30561 22457 30573 22460
rect 30607 22457 30619 22491
rect 30561 22451 30619 22457
rect 30834 22448 30840 22500
rect 30892 22488 30898 22500
rect 30892 22460 33548 22488
rect 30892 22448 30898 22460
rect 23808 22392 25268 22420
rect 23808 22380 23814 22392
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 25774 22380 25780 22432
rect 25832 22420 25838 22432
rect 26510 22420 26516 22432
rect 25832 22392 26516 22420
rect 25832 22380 25838 22392
rect 26510 22380 26516 22392
rect 26568 22380 26574 22432
rect 26602 22380 26608 22432
rect 26660 22380 26666 22432
rect 27798 22380 27804 22432
rect 27856 22380 27862 22432
rect 29178 22380 29184 22432
rect 29236 22420 29242 22432
rect 30098 22420 30104 22432
rect 29236 22392 30104 22420
rect 29236 22380 29242 22392
rect 30098 22380 30104 22392
rect 30156 22380 30162 22432
rect 30190 22380 30196 22432
rect 30248 22420 30254 22432
rect 31754 22420 31760 22432
rect 30248 22392 31760 22420
rect 30248 22380 30254 22392
rect 31754 22380 31760 22392
rect 31812 22420 31818 22432
rect 32030 22420 32036 22432
rect 31812 22392 32036 22420
rect 31812 22380 31818 22392
rect 32030 22380 32036 22392
rect 32088 22420 32094 22432
rect 33226 22420 33232 22432
rect 32088 22392 33232 22420
rect 32088 22380 32094 22392
rect 33226 22380 33232 22392
rect 33284 22380 33290 22432
rect 33520 22420 33548 22460
rect 33594 22448 33600 22500
rect 33652 22488 33658 22500
rect 33689 22491 33747 22497
rect 33689 22488 33701 22491
rect 33652 22460 33701 22488
rect 33652 22448 33658 22460
rect 33689 22457 33701 22460
rect 33735 22457 33747 22491
rect 33796 22488 33824 22516
rect 36832 22488 36860 22596
rect 37826 22516 37832 22568
rect 37884 22556 37890 22568
rect 37936 22565 37964 22596
rect 37921 22559 37979 22565
rect 37921 22556 37933 22559
rect 37884 22528 37933 22556
rect 37884 22516 37890 22528
rect 37921 22525 37933 22528
rect 37967 22525 37979 22559
rect 37921 22519 37979 22525
rect 38197 22559 38255 22565
rect 38197 22525 38209 22559
rect 38243 22556 38255 22559
rect 48682 22556 48688 22568
rect 38243 22528 48688 22556
rect 38243 22525 38255 22528
rect 38197 22519 38255 22525
rect 48682 22516 48688 22528
rect 48740 22516 48746 22568
rect 40497 22491 40555 22497
rect 40497 22488 40509 22491
rect 33796 22460 36860 22488
rect 39224 22460 40509 22488
rect 33689 22451 33747 22457
rect 35894 22420 35900 22432
rect 33520 22392 35900 22420
rect 35894 22380 35900 22392
rect 35952 22380 35958 22432
rect 36078 22380 36084 22432
rect 36136 22420 36142 22432
rect 36541 22423 36599 22429
rect 36541 22420 36553 22423
rect 36136 22392 36553 22420
rect 36136 22380 36142 22392
rect 36541 22389 36553 22392
rect 36587 22389 36599 22423
rect 36541 22383 36599 22389
rect 36906 22380 36912 22432
rect 36964 22380 36970 22432
rect 38378 22380 38384 22432
rect 38436 22420 38442 22432
rect 39224 22420 39252 22460
rect 40497 22457 40509 22460
rect 40543 22488 40555 22491
rect 40862 22488 40868 22500
rect 40543 22460 40868 22488
rect 40543 22457 40555 22460
rect 40497 22451 40555 22457
rect 40862 22448 40868 22460
rect 40920 22448 40926 22500
rect 38436 22392 39252 22420
rect 39669 22423 39727 22429
rect 38436 22380 38442 22392
rect 39669 22389 39681 22423
rect 39715 22420 39727 22423
rect 39758 22420 39764 22432
rect 39715 22392 39764 22420
rect 39715 22389 39727 22392
rect 39669 22383 39727 22389
rect 39758 22380 39764 22392
rect 39816 22380 39822 22432
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 6638 22216 6644 22228
rect 4120 22188 6644 22216
rect 4120 22176 4126 22188
rect 6638 22176 6644 22188
rect 6696 22176 6702 22228
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 11146 22216 11152 22228
rect 9824 22188 11152 22216
rect 9824 22176 9830 22188
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 16298 22216 16304 22228
rect 11388 22188 16304 22216
rect 11388 22176 11394 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 17392 22219 17450 22225
rect 17392 22185 17404 22219
rect 17438 22216 17450 22219
rect 17862 22216 17868 22228
rect 17438 22188 17868 22216
rect 17438 22185 17450 22188
rect 17392 22179 17450 22185
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 19334 22176 19340 22228
rect 19392 22216 19398 22228
rect 20073 22219 20131 22225
rect 20073 22216 20085 22219
rect 19392 22188 20085 22216
rect 19392 22176 19398 22188
rect 20073 22185 20085 22188
rect 20119 22216 20131 22219
rect 20438 22216 20444 22228
rect 20119 22188 20444 22216
rect 20119 22185 20131 22188
rect 20073 22179 20131 22185
rect 20438 22176 20444 22188
rect 20496 22176 20502 22228
rect 21450 22176 21456 22228
rect 21508 22216 21514 22228
rect 25130 22216 25136 22228
rect 21508 22188 25136 22216
rect 21508 22176 21514 22188
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 26040 22219 26098 22225
rect 26040 22185 26052 22219
rect 26086 22216 26098 22219
rect 27798 22216 27804 22228
rect 26086 22188 27804 22216
rect 26086 22185 26098 22188
rect 26040 22179 26098 22185
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 28902 22176 28908 22228
rect 28960 22216 28966 22228
rect 29273 22219 29331 22225
rect 29273 22216 29285 22219
rect 28960 22188 29285 22216
rect 28960 22176 28966 22188
rect 29273 22185 29285 22188
rect 29319 22216 29331 22219
rect 29549 22219 29607 22225
rect 29549 22216 29561 22219
rect 29319 22188 29561 22216
rect 29319 22185 29331 22188
rect 29273 22179 29331 22185
rect 29549 22185 29561 22188
rect 29595 22185 29607 22219
rect 31938 22216 31944 22228
rect 29549 22179 29607 22185
rect 29656 22188 31944 22216
rect 3786 22108 3792 22160
rect 3844 22148 3850 22160
rect 5534 22148 5540 22160
rect 3844 22120 5540 22148
rect 3844 22108 3850 22120
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 6104 22120 6592 22148
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3694 22040 3700 22092
rect 3752 22080 3758 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3752 22052 4445 22080
rect 3752 22040 3758 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 1780 21944 1808 21975
rect 4062 21972 4068 22024
rect 4120 21972 4126 22024
rect 6104 22012 6132 22120
rect 6564 22080 6592 22120
rect 6914 22108 6920 22160
rect 6972 22148 6978 22160
rect 10686 22148 10692 22160
rect 6972 22120 7328 22148
rect 6972 22108 6978 22120
rect 7300 22089 7328 22120
rect 9646 22120 10692 22148
rect 7285 22083 7343 22089
rect 6564 22052 6960 22080
rect 4356 21984 6132 22012
rect 6365 22015 6423 22021
rect 4154 21944 4160 21956
rect 1780 21916 4160 21944
rect 4154 21904 4160 21916
rect 4212 21904 4218 21956
rect 4356 21888 4384 21984
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 21981 6883 22015
rect 6932 22012 6960 22052
rect 7285 22049 7297 22083
rect 7331 22049 7343 22083
rect 7285 22043 7343 22049
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 7834 22080 7840 22092
rect 7616 22052 7840 22080
rect 7616 22040 7622 22052
rect 7834 22040 7840 22052
rect 7892 22040 7898 22092
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 9646 22080 9674 22120
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 10870 22108 10876 22160
rect 10928 22148 10934 22160
rect 10928 22120 13492 22148
rect 10928 22108 10934 22120
rect 8803 22052 9674 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 9950 22040 9956 22092
rect 10008 22040 10014 22092
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 11348 22052 12480 22080
rect 10502 22012 10508 22024
rect 6932 21984 10508 22012
rect 6825 21975 6883 21981
rect 5626 21904 5632 21956
rect 5684 21904 5690 21956
rect 3418 21836 3424 21888
rect 3476 21836 3482 21888
rect 3605 21879 3663 21885
rect 3605 21845 3617 21879
rect 3651 21876 3663 21879
rect 4338 21876 4344 21888
rect 3651 21848 4344 21876
rect 3651 21845 3663 21848
rect 3605 21839 3663 21845
rect 4338 21836 4344 21848
rect 4396 21836 4402 21888
rect 5902 21836 5908 21888
rect 5960 21836 5966 21888
rect 6178 21836 6184 21888
rect 6236 21836 6242 21888
rect 6380 21876 6408 21975
rect 6840 21944 6868 21975
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 10870 21972 10876 22024
rect 10928 22012 10934 22024
rect 11348 22012 11376 22052
rect 10928 21984 11376 22012
rect 10928 21972 10934 21984
rect 12342 21972 12348 22024
rect 12400 21972 12406 22024
rect 12452 22012 12480 22052
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 13464 22080 13492 22120
rect 13906 22108 13912 22160
rect 13964 22148 13970 22160
rect 14093 22151 14151 22157
rect 14093 22148 14105 22151
rect 13964 22120 14105 22148
rect 13964 22108 13970 22120
rect 14093 22117 14105 22120
rect 14139 22148 14151 22151
rect 14550 22148 14556 22160
rect 14139 22120 14556 22148
rect 14139 22117 14151 22120
rect 14093 22111 14151 22117
rect 14550 22108 14556 22120
rect 14608 22108 14614 22160
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 15160 22120 15700 22148
rect 15160 22108 15166 22120
rect 15672 22089 15700 22120
rect 20622 22108 20628 22160
rect 20680 22148 20686 22160
rect 21818 22148 21824 22160
rect 20680 22120 21824 22148
rect 20680 22108 20686 22120
rect 21818 22108 21824 22120
rect 21876 22108 21882 22160
rect 23290 22108 23296 22160
rect 23348 22108 23354 22160
rect 25774 22148 25780 22160
rect 23952 22120 25780 22148
rect 15657 22083 15715 22089
rect 13464 22052 15424 22080
rect 13078 22012 13084 22024
rect 12452 21984 13084 22012
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 15396 22021 15424 22052
rect 15657 22049 15669 22083
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 17129 22083 17187 22089
rect 17129 22049 17141 22083
rect 17175 22080 17187 22083
rect 19426 22080 19432 22092
rect 17175 22052 19432 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 19426 22040 19432 22052
rect 19484 22080 19490 22092
rect 19702 22080 19708 22092
rect 19484 22052 19708 22080
rect 19484 22040 19490 22052
rect 19702 22040 19708 22052
rect 19760 22040 19766 22092
rect 20530 22040 20536 22092
rect 20588 22080 20594 22092
rect 23952 22089 23980 22120
rect 25774 22108 25780 22120
rect 25832 22108 25838 22160
rect 27525 22151 27583 22157
rect 27525 22117 27537 22151
rect 27571 22148 27583 22151
rect 28350 22148 28356 22160
rect 27571 22120 28356 22148
rect 27571 22117 27583 22120
rect 27525 22111 27583 22117
rect 28350 22108 28356 22120
rect 28408 22148 28414 22160
rect 29656 22148 29684 22188
rect 31938 22176 31944 22188
rect 31996 22176 32002 22228
rect 32490 22176 32496 22228
rect 32548 22216 32554 22228
rect 36262 22216 36268 22228
rect 32548 22188 36268 22216
rect 32548 22176 32554 22188
rect 36262 22176 36268 22188
rect 36320 22176 36326 22228
rect 37553 22219 37611 22225
rect 37553 22185 37565 22219
rect 37599 22216 37611 22219
rect 38286 22216 38292 22228
rect 37599 22188 38292 22216
rect 37599 22185 37611 22188
rect 37553 22179 37611 22185
rect 38286 22176 38292 22188
rect 38344 22176 38350 22228
rect 39482 22216 39488 22228
rect 38396 22188 39488 22216
rect 28408 22120 29684 22148
rect 28408 22108 28414 22120
rect 30558 22108 30564 22160
rect 30616 22108 30622 22160
rect 31110 22108 31116 22160
rect 31168 22148 31174 22160
rect 34333 22151 34391 22157
rect 34333 22148 34345 22151
rect 31168 22120 34345 22148
rect 31168 22108 31174 22120
rect 34333 22117 34345 22120
rect 34379 22117 34391 22151
rect 34333 22111 34391 22117
rect 34422 22108 34428 22160
rect 34480 22148 34486 22160
rect 38396 22148 38424 22188
rect 39482 22176 39488 22188
rect 39540 22176 39546 22228
rect 34480 22120 38424 22148
rect 34480 22108 34486 22120
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 20588 22052 20821 22080
rect 20588 22040 20594 22052
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 24854 22080 24860 22092
rect 23983 22052 24017 22080
rect 24228 22052 24860 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 13188 21984 14565 22012
rect 7742 21944 7748 21956
rect 6840 21916 7748 21944
rect 7742 21904 7748 21916
rect 7800 21904 7806 21956
rect 8846 21944 8852 21956
rect 8220 21916 8852 21944
rect 8220 21876 8248 21916
rect 8846 21904 8852 21916
rect 8904 21904 8910 21956
rect 9033 21947 9091 21953
rect 9033 21913 9045 21947
rect 9079 21944 9091 21947
rect 9079 21916 10732 21944
rect 9079 21913 9091 21916
rect 9033 21907 9091 21913
rect 6380 21848 8248 21876
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 8481 21879 8539 21885
rect 8481 21876 8493 21879
rect 8352 21848 8493 21876
rect 8352 21836 8358 21848
rect 8481 21845 8493 21848
rect 8527 21845 8539 21879
rect 8864 21876 8892 21904
rect 9214 21876 9220 21888
rect 8864 21848 9220 21876
rect 8481 21839 8539 21845
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 10594 21876 10600 21888
rect 9723 21848 10600 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 10704 21876 10732 21916
rect 11054 21904 11060 21956
rect 11112 21944 11118 21956
rect 13188 21944 13216 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 15562 22012 15568 22024
rect 15427 21984 15568 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 18840 21984 20361 22012
rect 18840 21972 18846 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 22189 22015 22247 22021
rect 22189 21981 22201 22015
rect 22235 22012 22247 22015
rect 22646 22012 22652 22024
rect 22235 21984 22652 22012
rect 22235 21981 22247 21984
rect 22189 21975 22247 21981
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 23658 21972 23664 22024
rect 23716 21972 23722 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 24228 22012 24256 22052
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 25130 22040 25136 22092
rect 25188 22080 25194 22092
rect 25225 22083 25283 22089
rect 25225 22080 25237 22083
rect 25188 22052 25237 22080
rect 25188 22040 25194 22052
rect 25225 22049 25237 22052
rect 25271 22080 25283 22083
rect 25271 22052 29316 22080
rect 25271 22049 25283 22052
rect 25225 22043 25283 22049
rect 23799 21984 24256 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 24302 21972 24308 22024
rect 24360 22012 24366 22024
rect 25777 22015 25835 22021
rect 25777 22012 25789 22015
rect 24360 21984 25789 22012
rect 24360 21972 24366 21984
rect 25777 21981 25789 21984
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 27985 22015 28043 22021
rect 27985 22012 27997 22015
rect 27856 21984 27997 22012
rect 27856 21972 27862 21984
rect 27985 21981 27997 21984
rect 28031 21981 28043 22015
rect 27985 21975 28043 21981
rect 11112 21916 13216 21944
rect 11112 21904 11118 21916
rect 14090 21904 14096 21956
rect 14148 21944 14154 21956
rect 14148 21916 17816 21944
rect 14148 21904 14154 21916
rect 14274 21876 14280 21888
rect 10704 21848 14280 21876
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 14642 21836 14648 21888
rect 14700 21836 14706 21888
rect 14918 21836 14924 21888
rect 14976 21876 14982 21888
rect 15102 21876 15108 21888
rect 14976 21848 15108 21876
rect 14976 21836 14982 21848
rect 15102 21836 15108 21848
rect 15160 21876 15166 21888
rect 16114 21876 16120 21888
rect 15160 21848 16120 21876
rect 15160 21836 15166 21848
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 17788 21876 17816 21916
rect 17862 21904 17868 21956
rect 17920 21904 17926 21956
rect 19518 21944 19524 21956
rect 18708 21916 19524 21944
rect 18708 21876 18736 21916
rect 19518 21904 19524 21916
rect 19576 21904 19582 21956
rect 25041 21947 25099 21953
rect 22066 21916 24624 21944
rect 17788 21848 18736 21876
rect 18874 21836 18880 21888
rect 18932 21836 18938 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 19334 21876 19340 21888
rect 19300 21848 19340 21876
rect 19300 21836 19306 21848
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 19610 21836 19616 21888
rect 19668 21836 19674 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 22066 21876 22094 21916
rect 20128 21848 22094 21876
rect 22833 21879 22891 21885
rect 20128 21836 20134 21848
rect 22833 21845 22845 21879
rect 22879 21876 22891 21879
rect 24486 21876 24492 21888
rect 22879 21848 24492 21876
rect 22879 21845 22891 21848
rect 22833 21839 22891 21845
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24596 21885 24624 21916
rect 25041 21913 25053 21947
rect 25087 21944 25099 21947
rect 25498 21944 25504 21956
rect 25087 21916 25504 21944
rect 25087 21913 25099 21916
rect 25041 21907 25099 21913
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 25590 21904 25596 21956
rect 25648 21944 25654 21956
rect 26050 21944 26056 21956
rect 25648 21916 26056 21944
rect 25648 21904 25654 21916
rect 26050 21904 26056 21916
rect 26108 21944 26114 21956
rect 26510 21944 26516 21956
rect 26108 21916 26516 21944
rect 26108 21904 26114 21916
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 29178 21944 29184 21956
rect 27396 21916 29184 21944
rect 27396 21904 27402 21916
rect 29178 21904 29184 21916
rect 29236 21904 29242 21956
rect 29288 21944 29316 22052
rect 29362 22040 29368 22092
rect 29420 22080 29426 22092
rect 30282 22080 30288 22092
rect 29420 22052 30288 22080
rect 29420 22040 29426 22052
rect 30282 22040 30288 22052
rect 30340 22040 30346 22092
rect 30469 22083 30527 22089
rect 30469 22049 30481 22083
rect 30515 22080 30527 22083
rect 30576 22080 30604 22108
rect 30515 22052 30604 22080
rect 30515 22049 30527 22052
rect 30469 22043 30527 22049
rect 30650 22040 30656 22092
rect 30708 22040 30714 22092
rect 31018 22040 31024 22092
rect 31076 22080 31082 22092
rect 31076 22052 32720 22080
rect 31076 22040 31082 22052
rect 30098 21972 30104 22024
rect 30156 22012 30162 22024
rect 31205 22015 31263 22021
rect 31205 22012 31217 22015
rect 30156 21984 31217 22012
rect 30156 21972 30162 21984
rect 31205 21981 31217 21984
rect 31251 21981 31263 22015
rect 32309 22015 32367 22021
rect 32309 22012 32321 22015
rect 31205 21975 31263 21981
rect 31726 21984 32321 22012
rect 31726 21944 31754 21984
rect 32309 21981 32321 21984
rect 32355 21981 32367 22015
rect 32692 22012 32720 22052
rect 32766 22040 32772 22092
rect 32824 22080 32830 22092
rect 32953 22083 33011 22089
rect 32953 22080 32965 22083
rect 32824 22052 32965 22080
rect 32824 22040 32830 22052
rect 32953 22049 32965 22052
rect 32999 22049 33011 22083
rect 35161 22083 35219 22089
rect 32953 22043 33011 22049
rect 33060 22052 35112 22080
rect 33060 22012 33088 22052
rect 32692 21984 33088 22012
rect 33413 22015 33471 22021
rect 32309 21975 32367 21981
rect 33413 21981 33425 22015
rect 33459 21981 33471 22015
rect 35084 22012 35112 22052
rect 35161 22049 35173 22083
rect 35207 22080 35219 22083
rect 35250 22080 35256 22092
rect 35207 22052 35256 22080
rect 35207 22049 35219 22052
rect 35161 22043 35219 22049
rect 35250 22040 35256 22052
rect 35308 22040 35314 22092
rect 36262 22040 36268 22092
rect 36320 22080 36326 22092
rect 39669 22083 39727 22089
rect 36320 22052 39068 22080
rect 36320 22040 36326 22052
rect 35084 21984 37044 22012
rect 33413 21975 33471 21981
rect 29288 21916 31754 21944
rect 31938 21904 31944 21956
rect 31996 21944 32002 21956
rect 33428 21944 33456 21975
rect 31996 21916 33456 21944
rect 31996 21904 32002 21916
rect 33870 21904 33876 21956
rect 33928 21944 33934 21956
rect 33928 21916 34192 21944
rect 33928 21904 33934 21916
rect 24581 21879 24639 21885
rect 24581 21845 24593 21879
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 24946 21836 24952 21888
rect 25004 21836 25010 21888
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 26292 21848 28641 21876
rect 26292 21836 26298 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 28997 21879 29055 21885
rect 28997 21845 29009 21879
rect 29043 21876 29055 21879
rect 29086 21876 29092 21888
rect 29043 21848 29092 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29086 21836 29092 21848
rect 29144 21876 29150 21888
rect 29362 21876 29368 21888
rect 29144 21848 29368 21876
rect 29144 21836 29150 21848
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 30006 21836 30012 21888
rect 30064 21836 30070 21888
rect 30282 21836 30288 21888
rect 30340 21876 30346 21888
rect 30377 21879 30435 21885
rect 30377 21876 30389 21879
rect 30340 21848 30389 21876
rect 30340 21836 30346 21848
rect 30377 21845 30389 21848
rect 30423 21845 30435 21879
rect 30377 21839 30435 21845
rect 30466 21836 30472 21888
rect 30524 21876 30530 21888
rect 31849 21879 31907 21885
rect 31849 21876 31861 21879
rect 30524 21848 31861 21876
rect 30524 21836 30530 21848
rect 31849 21845 31861 21848
rect 31895 21845 31907 21879
rect 31849 21839 31907 21845
rect 32122 21836 32128 21888
rect 32180 21876 32186 21888
rect 34057 21879 34115 21885
rect 34057 21876 34069 21879
rect 32180 21848 34069 21876
rect 32180 21836 32186 21848
rect 34057 21845 34069 21848
rect 34103 21845 34115 21879
rect 34164 21876 34192 21916
rect 34606 21904 34612 21956
rect 34664 21944 34670 21956
rect 34977 21947 35035 21953
rect 34977 21944 34989 21947
rect 34664 21916 34989 21944
rect 34664 21904 34670 21916
rect 34977 21913 34989 21916
rect 35023 21913 35035 21947
rect 34977 21907 35035 21913
rect 35710 21904 35716 21956
rect 35768 21904 35774 21956
rect 35894 21904 35900 21956
rect 35952 21904 35958 21956
rect 36909 21947 36967 21953
rect 36909 21913 36921 21947
rect 36955 21913 36967 21947
rect 37016 21944 37044 21984
rect 37090 21972 37096 22024
rect 37148 21972 37154 22024
rect 37734 21972 37740 22024
rect 37792 21972 37798 22024
rect 37918 21972 37924 22024
rect 37976 22012 37982 22024
rect 38286 22012 38292 22024
rect 37976 21984 38292 22012
rect 37976 21972 37982 21984
rect 38286 21972 38292 21984
rect 38344 22012 38350 22024
rect 39040 22021 39068 22052
rect 39669 22049 39681 22083
rect 39715 22080 39727 22083
rect 39850 22080 39856 22092
rect 39715 22052 39856 22080
rect 39715 22049 39727 22052
rect 39669 22043 39727 22049
rect 39850 22040 39856 22052
rect 39908 22040 39914 22092
rect 38381 22015 38439 22021
rect 38381 22012 38393 22015
rect 38344 21984 38393 22012
rect 38344 21972 38350 21984
rect 38381 21981 38393 21984
rect 38427 21981 38439 22015
rect 38381 21975 38439 21981
rect 39025 22015 39083 22021
rect 39025 21981 39037 22015
rect 39071 22012 39083 22015
rect 39301 22015 39359 22021
rect 39301 22012 39313 22015
rect 39071 21984 39313 22012
rect 39071 21981 39083 21984
rect 39025 21975 39083 21981
rect 39301 21981 39313 21984
rect 39347 21981 39359 22015
rect 39301 21975 39359 21981
rect 37016 21916 38654 21944
rect 36909 21907 36967 21913
rect 36173 21879 36231 21885
rect 36173 21876 36185 21879
rect 34164 21848 36185 21876
rect 34057 21839 34115 21845
rect 36173 21845 36185 21848
rect 36219 21845 36231 21879
rect 36173 21839 36231 21845
rect 36262 21836 36268 21888
rect 36320 21876 36326 21888
rect 36357 21879 36415 21885
rect 36357 21876 36369 21879
rect 36320 21848 36369 21876
rect 36320 21836 36326 21848
rect 36357 21845 36369 21848
rect 36403 21845 36415 21879
rect 36924 21876 36952 21907
rect 37090 21876 37096 21888
rect 36924 21848 37096 21876
rect 36357 21839 36415 21845
rect 37090 21836 37096 21848
rect 37148 21836 37154 21888
rect 37182 21836 37188 21888
rect 37240 21876 37246 21888
rect 38197 21879 38255 21885
rect 38197 21876 38209 21879
rect 37240 21848 38209 21876
rect 37240 21836 37246 21848
rect 38197 21845 38209 21848
rect 38243 21845 38255 21879
rect 38626 21876 38654 21916
rect 38841 21879 38899 21885
rect 38841 21876 38853 21879
rect 38626 21848 38853 21876
rect 38197 21839 38255 21845
rect 38841 21845 38853 21848
rect 38887 21845 38899 21879
rect 38841 21839 38899 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 6914 21672 6920 21684
rect 4212 21644 6920 21672
rect 4212 21632 4218 21644
rect 6914 21632 6920 21644
rect 6972 21632 6978 21684
rect 7101 21675 7159 21681
rect 7101 21641 7113 21675
rect 7147 21672 7159 21675
rect 8478 21672 8484 21684
rect 7147 21644 8484 21672
rect 7147 21641 7159 21644
rect 7101 21635 7159 21641
rect 8478 21632 8484 21644
rect 8536 21632 8542 21684
rect 9585 21675 9643 21681
rect 9585 21641 9597 21675
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 10870 21672 10876 21684
rect 10183 21644 10876 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 3234 21604 3240 21616
rect 1780 21576 3240 21604
rect 1780 21545 1808 21576
rect 3234 21564 3240 21576
rect 3292 21564 3298 21616
rect 3694 21564 3700 21616
rect 3752 21604 3758 21616
rect 5721 21607 5779 21613
rect 5721 21604 5733 21607
rect 3752 21576 5733 21604
rect 3752 21564 3758 21576
rect 5721 21573 5733 21576
rect 5767 21573 5779 21607
rect 5721 21567 5779 21573
rect 6656 21576 7788 21604
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21505 1823 21539
rect 1765 21499 1823 21505
rect 2314 21496 2320 21548
rect 2372 21536 2378 21548
rect 3421 21539 3479 21545
rect 3421 21536 3433 21539
rect 2372 21508 3433 21536
rect 2372 21496 2378 21508
rect 3421 21505 3433 21508
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 6656 21536 6684 21576
rect 7009 21539 7067 21545
rect 7009 21536 7021 21539
rect 5675 21508 6684 21536
rect 6748 21508 7021 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3326 21468 3332 21480
rect 2823 21440 3332 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 3881 21471 3939 21477
rect 3881 21468 3893 21471
rect 3660 21440 3893 21468
rect 3660 21428 3666 21440
rect 3881 21437 3893 21440
rect 3927 21437 3939 21471
rect 3881 21431 3939 21437
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6086 21468 6092 21480
rect 5951 21440 6092 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 1118 21360 1124 21412
rect 1176 21400 1182 21412
rect 6641 21403 6699 21409
rect 6641 21400 6653 21403
rect 1176 21372 6653 21400
rect 1176 21360 1182 21372
rect 6641 21369 6653 21372
rect 6687 21369 6699 21403
rect 6641 21363 6699 21369
rect 3234 21292 3240 21344
rect 3292 21332 3298 21344
rect 3418 21332 3424 21344
rect 3292 21304 3424 21332
rect 3292 21292 3298 21304
rect 3418 21292 3424 21304
rect 3476 21292 3482 21344
rect 4982 21292 4988 21344
rect 5040 21332 5046 21344
rect 5261 21335 5319 21341
rect 5261 21332 5273 21335
rect 5040 21304 5273 21332
rect 5040 21292 5046 21304
rect 5261 21301 5273 21304
rect 5307 21301 5319 21335
rect 5261 21295 5319 21301
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 6457 21335 6515 21341
rect 6457 21332 6469 21335
rect 5500 21304 6469 21332
rect 5500 21292 5506 21304
rect 6457 21301 6469 21304
rect 6503 21332 6515 21335
rect 6748 21332 6776 21508
rect 7009 21505 7021 21508
rect 7055 21536 7067 21539
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 7055 21508 7481 21536
rect 7055 21505 7067 21508
rect 7009 21499 7067 21505
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7190 21428 7196 21480
rect 7248 21428 7254 21480
rect 7098 21360 7104 21412
rect 7156 21400 7162 21412
rect 7558 21400 7564 21412
rect 7156 21372 7564 21400
rect 7156 21360 7162 21372
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 7760 21400 7788 21576
rect 8110 21564 8116 21616
rect 8168 21564 8174 21616
rect 9122 21564 9128 21616
rect 9180 21564 9186 21616
rect 9600 21604 9628 21635
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 10962 21632 10968 21684
rect 11020 21672 11026 21684
rect 11977 21675 12035 21681
rect 11977 21672 11989 21675
rect 11020 21644 11989 21672
rect 11020 21632 11026 21644
rect 11977 21641 11989 21644
rect 12023 21641 12035 21675
rect 11977 21635 12035 21641
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 12492 21644 13216 21672
rect 12492 21632 12498 21644
rect 11790 21604 11796 21616
rect 9600 21576 11796 21604
rect 11790 21564 11796 21576
rect 11848 21604 11854 21616
rect 12526 21604 12532 21616
rect 11848 21576 12532 21604
rect 11848 21564 11854 21576
rect 12526 21564 12532 21576
rect 12584 21564 12590 21616
rect 13188 21604 13216 21644
rect 14274 21632 14280 21684
rect 14332 21672 14338 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 14332 21644 15945 21672
rect 14332 21632 14338 21644
rect 15933 21641 15945 21644
rect 15979 21672 15991 21675
rect 17773 21675 17831 21681
rect 17773 21672 17785 21675
rect 15979 21644 17785 21672
rect 15979 21641 15991 21644
rect 15933 21635 15991 21641
rect 17773 21641 17785 21644
rect 17819 21672 17831 21675
rect 22465 21675 22523 21681
rect 17819 21644 22094 21672
rect 17819 21641 17831 21644
rect 17773 21635 17831 21641
rect 13722 21604 13728 21616
rect 13188 21576 13728 21604
rect 9766 21496 9772 21548
rect 9824 21536 9830 21548
rect 10781 21539 10839 21545
rect 10781 21536 10793 21539
rect 9824 21508 10793 21536
rect 9824 21496 9830 21508
rect 10781 21505 10793 21508
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 11664 21508 12357 21536
rect 11664 21496 11670 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 7834 21428 7840 21480
rect 7892 21428 7898 21480
rect 10318 21468 10324 21480
rect 7944 21440 10324 21468
rect 7944 21400 7972 21440
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10870 21428 10876 21480
rect 10928 21428 10934 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 12544 21477 12572 21564
rect 13188 21545 13216 21576
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 14918 21564 14924 21616
rect 14976 21604 14982 21616
rect 18782 21604 18788 21616
rect 14976 21576 18788 21604
rect 14976 21564 14982 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 19334 21564 19340 21616
rect 19392 21564 19398 21616
rect 22066 21604 22094 21644
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22511 21644 24992 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23198 21604 23204 21616
rect 22066 21576 23204 21604
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 23661 21607 23719 21613
rect 23661 21604 23673 21607
rect 23624 21576 23673 21604
rect 23624 21564 23630 21576
rect 23661 21573 23673 21576
rect 23707 21573 23719 21607
rect 23661 21567 23719 21573
rect 23934 21564 23940 21616
rect 23992 21604 23998 21616
rect 24964 21604 24992 21644
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 25961 21675 26019 21681
rect 25961 21672 25973 21675
rect 25096 21644 25973 21672
rect 25096 21632 25102 21644
rect 25961 21641 25973 21644
rect 26007 21641 26019 21675
rect 25961 21635 26019 21641
rect 26142 21632 26148 21684
rect 26200 21672 26206 21684
rect 27249 21675 27307 21681
rect 27249 21672 27261 21675
rect 26200 21644 27261 21672
rect 26200 21632 26206 21644
rect 27249 21641 27261 21644
rect 27295 21641 27307 21675
rect 27249 21635 27307 21641
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 28626 21672 28632 21684
rect 27755 21644 28632 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 28626 21632 28632 21644
rect 28684 21632 28690 21684
rect 30006 21672 30012 21684
rect 29104 21644 30012 21672
rect 25314 21604 25320 21616
rect 23992 21576 24150 21604
rect 24964 21576 25320 21604
rect 23992 21564 23998 21576
rect 25314 21564 25320 21576
rect 25372 21564 25378 21616
rect 26053 21607 26111 21613
rect 26053 21573 26065 21607
rect 26099 21604 26111 21607
rect 29104 21604 29132 21644
rect 30006 21632 30012 21644
rect 30064 21632 30070 21684
rect 30650 21632 30656 21684
rect 30708 21632 30714 21684
rect 31018 21632 31024 21684
rect 31076 21632 31082 21684
rect 31113 21675 31171 21681
rect 31113 21641 31125 21675
rect 31159 21672 31171 21675
rect 33226 21672 33232 21684
rect 31159 21644 33232 21672
rect 31159 21641 31171 21644
rect 31113 21635 31171 21641
rect 33226 21632 33232 21644
rect 33284 21632 33290 21684
rect 33410 21632 33416 21684
rect 33468 21632 33474 21684
rect 34698 21632 34704 21684
rect 34756 21632 34762 21684
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 35989 21675 36047 21681
rect 35989 21672 36001 21675
rect 35943 21644 36001 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 35989 21641 36001 21644
rect 36035 21672 36047 21675
rect 36170 21672 36176 21684
rect 36035 21644 36176 21672
rect 36035 21641 36047 21644
rect 35989 21635 36047 21641
rect 36170 21632 36176 21644
rect 36228 21632 36234 21684
rect 36814 21632 36820 21684
rect 36872 21672 36878 21684
rect 37461 21675 37519 21681
rect 37461 21672 37473 21675
rect 36872 21644 37473 21672
rect 36872 21632 36878 21644
rect 37461 21641 37473 21644
rect 37507 21641 37519 21675
rect 37461 21635 37519 21641
rect 37826 21632 37832 21684
rect 37884 21672 37890 21684
rect 38381 21675 38439 21681
rect 38381 21672 38393 21675
rect 37884 21644 38393 21672
rect 37884 21632 37890 21644
rect 38381 21641 38393 21644
rect 38427 21641 38439 21675
rect 38381 21635 38439 21641
rect 26099 21576 29132 21604
rect 26099 21573 26111 21576
rect 26053 21567 26111 21573
rect 29362 21564 29368 21616
rect 29420 21564 29426 21616
rect 30742 21564 30748 21616
rect 30800 21604 30806 21616
rect 34057 21607 34115 21613
rect 34057 21604 34069 21607
rect 30800 21576 34069 21604
rect 30800 21564 30806 21576
rect 34057 21573 34069 21576
rect 34103 21573 34115 21607
rect 34057 21567 34115 21573
rect 34330 21564 34336 21616
rect 34388 21604 34394 21616
rect 34388 21576 35480 21604
rect 34388 21564 34394 21576
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21505 13231 21539
rect 13173 21499 13231 21505
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 15197 21539 15255 21545
rect 15197 21536 15209 21539
rect 14608 21508 15209 21536
rect 14608 21496 14614 21508
rect 15197 21505 15209 21508
rect 15243 21536 15255 21539
rect 16666 21536 16672 21548
rect 15243 21508 16672 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 16666 21496 16672 21508
rect 16724 21536 16730 21548
rect 17770 21536 17776 21548
rect 16724 21508 17776 21536
rect 16724 21496 16730 21508
rect 17770 21496 17776 21508
rect 17828 21536 17834 21548
rect 18506 21536 18512 21548
rect 17828 21508 18512 21536
rect 17828 21496 17834 21508
rect 18506 21496 18512 21508
rect 18564 21496 18570 21548
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 20956 21508 22385 21536
rect 20956 21496 20962 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 25038 21496 25044 21548
rect 25096 21536 25102 21548
rect 27246 21536 27252 21548
rect 25096 21508 27252 21536
rect 25096 21496 25102 21508
rect 27246 21496 27252 21508
rect 27304 21536 27310 21548
rect 27522 21536 27528 21548
rect 27304 21508 27528 21536
rect 27304 21496 27310 21508
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21536 27675 21539
rect 27706 21536 27712 21548
rect 27663 21508 27712 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 27706 21496 27712 21508
rect 27764 21536 27770 21548
rect 28350 21536 28356 21548
rect 27764 21508 28356 21536
rect 27764 21496 27770 21508
rect 28350 21496 28356 21508
rect 28408 21496 28414 21548
rect 30282 21496 30288 21548
rect 30340 21536 30346 21548
rect 31757 21539 31815 21545
rect 31757 21536 31769 21539
rect 30340 21508 31769 21536
rect 30340 21496 30346 21508
rect 31757 21505 31769 21508
rect 31803 21536 31815 21539
rect 32214 21536 32220 21548
rect 31803 21508 32220 21536
rect 31803 21505 31815 21508
rect 31757 21499 31815 21505
rect 32214 21496 32220 21508
rect 32272 21496 32278 21548
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 34609 21539 34667 21545
rect 32824 21508 34008 21536
rect 32824 21496 32830 21508
rect 12437 21471 12495 21477
rect 12437 21468 12449 21471
rect 12216 21440 12449 21468
rect 12216 21428 12222 21440
rect 12437 21437 12449 21440
rect 12483 21437 12495 21471
rect 12437 21431 12495 21437
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21437 12587 21471
rect 12529 21431 12587 21437
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 12860 21440 13461 21468
rect 12860 21428 12866 21440
rect 13449 21437 13461 21440
rect 13495 21468 13507 21471
rect 13538 21468 13544 21480
rect 13495 21440 13544 21468
rect 13495 21437 13507 21440
rect 13449 21431 13507 21437
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 14921 21471 14979 21477
rect 14921 21468 14933 21471
rect 14056 21440 14933 21468
rect 14056 21428 14062 21440
rect 14921 21437 14933 21440
rect 14967 21437 14979 21471
rect 14921 21431 14979 21437
rect 16022 21428 16028 21480
rect 16080 21428 16086 21480
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21437 16175 21471
rect 16117 21431 16175 21437
rect 10778 21400 10784 21412
rect 7760 21372 7972 21400
rect 9140 21372 10784 21400
rect 6503 21304 6776 21332
rect 6503 21301 6515 21304
rect 6457 21295 6515 21301
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 9140 21332 9168 21372
rect 10778 21360 10784 21372
rect 10836 21360 10842 21412
rect 11514 21360 11520 21412
rect 11572 21400 11578 21412
rect 12710 21400 12716 21412
rect 11572 21372 12716 21400
rect 11572 21360 11578 21372
rect 12710 21360 12716 21372
rect 12768 21360 12774 21412
rect 16132 21400 16160 21431
rect 16942 21428 16948 21480
rect 17000 21428 17006 21480
rect 17126 21428 17132 21480
rect 17184 21468 17190 21480
rect 17862 21468 17868 21480
rect 17184 21440 17868 21468
rect 17184 21428 17190 21440
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 17957 21471 18015 21477
rect 17957 21437 17969 21471
rect 18003 21437 18015 21471
rect 17957 21431 18015 21437
rect 17678 21400 17684 21412
rect 15488 21372 17684 21400
rect 6972 21304 9168 21332
rect 6972 21292 6978 21304
rect 10410 21292 10416 21344
rect 10468 21292 10474 21344
rect 11422 21292 11428 21344
rect 11480 21332 11486 21344
rect 11609 21335 11667 21341
rect 11609 21332 11621 21335
rect 11480 21304 11621 21332
rect 11480 21292 11486 21304
rect 11609 21301 11621 21304
rect 11655 21301 11667 21335
rect 11609 21295 11667 21301
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 15488 21332 15516 21372
rect 17678 21360 17684 21372
rect 17736 21360 17742 21412
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 17972 21400 18000 21431
rect 18598 21428 18604 21480
rect 18656 21428 18662 21480
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 22704 21440 25145 21468
rect 22704 21428 22710 21440
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 26145 21471 26203 21477
rect 26145 21437 26157 21471
rect 26191 21468 26203 21471
rect 27338 21468 27344 21480
rect 26191 21440 27344 21468
rect 26191 21437 26203 21440
rect 26145 21431 26203 21437
rect 27338 21428 27344 21440
rect 27396 21428 27402 21480
rect 27798 21428 27804 21480
rect 27856 21428 27862 21480
rect 28445 21471 28503 21477
rect 28445 21437 28457 21471
rect 28491 21437 28503 21471
rect 28445 21431 28503 21437
rect 28721 21471 28779 21477
rect 28721 21437 28733 21471
rect 28767 21468 28779 21471
rect 30466 21468 30472 21480
rect 28767 21440 30472 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 22278 21400 22284 21412
rect 17828 21372 18000 21400
rect 20272 21372 22284 21400
rect 17828 21360 17834 21372
rect 13596 21304 15516 21332
rect 13596 21292 13602 21304
rect 15562 21292 15568 21344
rect 15620 21292 15626 21344
rect 17129 21335 17187 21341
rect 17129 21301 17141 21335
rect 17175 21332 17187 21335
rect 17218 21332 17224 21344
rect 17175 21304 17224 21332
rect 17175 21301 17187 21304
rect 17129 21295 17187 21301
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 17402 21292 17408 21344
rect 17460 21292 17466 21344
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 20272 21332 20300 21372
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 22370 21360 22376 21412
rect 22428 21400 22434 21412
rect 22428 21372 23520 21400
rect 22428 21360 22434 21372
rect 17552 21304 20300 21332
rect 20349 21335 20407 21341
rect 17552 21292 17558 21304
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20714 21332 20720 21344
rect 20395 21304 20720 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20714 21292 20720 21304
rect 20772 21292 20778 21344
rect 21450 21292 21456 21344
rect 21508 21292 21514 21344
rect 21542 21292 21548 21344
rect 21600 21332 21606 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21600 21304 22017 21332
rect 21600 21292 21606 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22005 21295 22063 21301
rect 23109 21335 23167 21341
rect 23109 21301 23121 21335
rect 23155 21332 23167 21335
rect 23382 21332 23388 21344
rect 23155 21304 23388 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23492 21332 23520 21372
rect 26694 21360 26700 21412
rect 26752 21400 26758 21412
rect 28460 21400 28488 21431
rect 30466 21428 30472 21440
rect 30524 21428 30530 21480
rect 31205 21471 31263 21477
rect 31205 21437 31217 21471
rect 31251 21437 31263 21471
rect 33873 21471 33931 21477
rect 33873 21468 33885 21471
rect 31205 21431 31263 21437
rect 31726 21440 33885 21468
rect 26752 21372 28488 21400
rect 26752 21360 26758 21372
rect 25593 21335 25651 21341
rect 25593 21332 25605 21335
rect 23492 21304 25605 21332
rect 25593 21301 25605 21304
rect 25639 21301 25651 21335
rect 25593 21295 25651 21301
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 26970 21332 26976 21344
rect 26016 21304 26976 21332
rect 26016 21292 26022 21304
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 28460 21332 28488 21372
rect 30193 21403 30251 21409
rect 30193 21369 30205 21403
rect 30239 21400 30251 21403
rect 30834 21400 30840 21412
rect 30239 21372 30840 21400
rect 30239 21369 30251 21372
rect 30193 21363 30251 21369
rect 30834 21360 30840 21372
rect 30892 21400 30898 21412
rect 31220 21400 31248 21431
rect 30892 21372 31248 21400
rect 30892 21360 30898 21372
rect 28902 21332 28908 21344
rect 28460 21304 28908 21332
rect 28902 21292 28908 21304
rect 28960 21292 28966 21344
rect 29086 21292 29092 21344
rect 29144 21332 29150 21344
rect 31018 21332 31024 21344
rect 29144 21304 31024 21332
rect 29144 21292 29150 21304
rect 31018 21292 31024 21304
rect 31076 21332 31082 21344
rect 31726 21332 31754 21440
rect 33873 21437 33885 21440
rect 33919 21437 33931 21471
rect 33980 21468 34008 21508
rect 34609 21505 34621 21539
rect 34655 21536 34667 21539
rect 34882 21536 34888 21548
rect 34655 21508 34888 21536
rect 34655 21505 34667 21508
rect 34609 21499 34667 21505
rect 34882 21496 34888 21508
rect 34940 21496 34946 21548
rect 35342 21496 35348 21548
rect 35400 21496 35406 21548
rect 35452 21536 35480 21576
rect 35526 21564 35532 21616
rect 35584 21604 35590 21616
rect 37277 21607 37335 21613
rect 37277 21604 37289 21607
rect 35584 21576 37289 21604
rect 35584 21564 35590 21576
rect 37277 21573 37289 21576
rect 37323 21573 37335 21607
rect 37277 21567 37335 21573
rect 38286 21564 38292 21616
rect 38344 21564 38350 21616
rect 36262 21536 36268 21548
rect 35452 21508 36268 21536
rect 36262 21496 36268 21508
rect 36320 21496 36326 21548
rect 36354 21496 36360 21548
rect 36412 21536 36418 21548
rect 36817 21539 36875 21545
rect 36817 21536 36829 21539
rect 36412 21508 36829 21536
rect 36412 21496 36418 21508
rect 36817 21505 36829 21508
rect 36863 21536 36875 21539
rect 37829 21539 37887 21545
rect 37829 21536 37841 21539
rect 36863 21508 37841 21536
rect 36863 21505 36875 21508
rect 36817 21499 36875 21505
rect 37829 21505 37841 21508
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 47578 21496 47584 21548
rect 47636 21536 47642 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47636 21508 47961 21536
rect 47636 21496 47642 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 35529 21471 35587 21477
rect 35529 21468 35541 21471
rect 33980 21440 35541 21468
rect 33873 21431 33931 21437
rect 35529 21437 35541 21440
rect 35575 21437 35587 21471
rect 35529 21431 35587 21437
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 31941 21403 31999 21409
rect 31941 21369 31953 21403
rect 31987 21400 31999 21403
rect 32030 21400 32036 21412
rect 31987 21372 32036 21400
rect 31987 21369 31999 21372
rect 31941 21363 31999 21369
rect 32030 21360 32036 21372
rect 32088 21360 32094 21412
rect 32214 21360 32220 21412
rect 32272 21400 32278 21412
rect 32272 21372 33180 21400
rect 32272 21360 32278 21372
rect 31076 21304 31754 21332
rect 31076 21292 31082 21304
rect 32122 21292 32128 21344
rect 32180 21332 32186 21344
rect 32953 21335 33011 21341
rect 32953 21332 32965 21335
rect 32180 21304 32965 21332
rect 32180 21292 32186 21304
rect 32953 21301 32965 21304
rect 32999 21301 33011 21335
rect 33152 21332 33180 21372
rect 33226 21360 33232 21412
rect 33284 21400 33290 21412
rect 36633 21403 36691 21409
rect 36633 21400 36645 21403
rect 33284 21372 36645 21400
rect 33284 21360 33290 21372
rect 36633 21369 36645 21372
rect 36679 21369 36691 21403
rect 36633 21363 36691 21369
rect 36722 21360 36728 21412
rect 36780 21400 36786 21412
rect 37645 21403 37703 21409
rect 37645 21400 37657 21403
rect 36780 21372 37657 21400
rect 36780 21360 36786 21372
rect 37645 21369 37657 21372
rect 37691 21369 37703 21403
rect 37645 21363 37703 21369
rect 34606 21332 34612 21344
rect 33152 21304 34612 21332
rect 32953 21295 33011 21301
rect 34606 21292 34612 21304
rect 34664 21332 34670 21344
rect 36906 21332 36912 21344
rect 34664 21304 36912 21332
rect 34664 21292 34670 21304
rect 36906 21292 36912 21304
rect 36964 21292 36970 21344
rect 37826 21292 37832 21344
rect 37884 21332 37890 21344
rect 38013 21335 38071 21341
rect 38013 21332 38025 21335
rect 37884 21304 38025 21332
rect 37884 21292 37890 21304
rect 38013 21301 38025 21304
rect 38059 21301 38071 21335
rect 38013 21295 38071 21301
rect 47578 21292 47584 21344
rect 47636 21292 47642 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3786 21088 3792 21140
rect 3844 21128 3850 21140
rect 3970 21128 3976 21140
rect 3844 21100 3976 21128
rect 3844 21088 3850 21100
rect 3970 21088 3976 21100
rect 4028 21088 4034 21140
rect 5810 21088 5816 21140
rect 5868 21088 5874 21140
rect 5902 21088 5908 21140
rect 5960 21128 5966 21140
rect 5960 21100 7604 21128
rect 5960 21088 5966 21100
rect 3421 21063 3479 21069
rect 3421 21029 3433 21063
rect 3467 21060 3479 21063
rect 5994 21060 6000 21072
rect 3467 21032 6000 21060
rect 3467 21029 3479 21032
rect 3421 21023 3479 21029
rect 5994 21020 6000 21032
rect 6052 21020 6058 21072
rect 7576 21060 7604 21100
rect 8018 21088 8024 21140
rect 8076 21088 8082 21140
rect 16022 21128 16028 21140
rect 8128 21100 16028 21128
rect 8128 21060 8156 21100
rect 16022 21088 16028 21100
rect 16080 21088 16086 21140
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 19061 21131 19119 21137
rect 16172 21100 17724 21128
rect 16172 21088 16178 21100
rect 7576 21032 8156 21060
rect 8757 21063 8815 21069
rect 8757 21029 8769 21063
rect 8803 21060 8815 21063
rect 13538 21060 13544 21072
rect 8803 21032 13544 21060
rect 8803 21029 8815 21032
rect 8757 21023 8815 21029
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 13725 21063 13783 21069
rect 13725 21029 13737 21063
rect 13771 21060 13783 21063
rect 13906 21060 13912 21072
rect 13771 21032 13912 21060
rect 13771 21029 13783 21032
rect 13725 21023 13783 21029
rect 13906 21020 13912 21032
rect 13964 21020 13970 21072
rect 17402 21060 17408 21072
rect 14200 21032 15424 21060
rect 3510 20952 3516 21004
rect 3568 20992 3574 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 3568 20964 4445 20992
rect 3568 20952 3574 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 6273 20995 6331 21001
rect 6273 20961 6285 20995
rect 6319 20992 6331 20995
rect 7834 20992 7840 21004
rect 6319 20964 7840 20992
rect 6319 20961 6331 20964
rect 6273 20955 6331 20961
rect 7834 20952 7840 20964
rect 7892 20952 7898 21004
rect 7926 20952 7932 21004
rect 7984 20992 7990 21004
rect 8297 20995 8355 21001
rect 8297 20992 8309 20995
rect 7984 20964 8309 20992
rect 7984 20952 7990 20964
rect 8297 20961 8309 20964
rect 8343 20992 8355 20995
rect 11514 20992 11520 21004
rect 8343 20964 11520 20992
rect 8343 20961 8355 20964
rect 8297 20955 8355 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 11882 20952 11888 21004
rect 11940 20992 11946 21004
rect 12437 20995 12495 21001
rect 12437 20992 12449 20995
rect 11940 20964 12449 20992
rect 11940 20952 11946 20964
rect 12437 20961 12449 20964
rect 12483 20961 12495 20995
rect 13446 20992 13452 21004
rect 12437 20955 12495 20961
rect 12636 20964 13452 20992
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1811 20896 3924 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 2866 20856 2872 20868
rect 2823 20828 2872 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 3896 20856 3924 20896
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 9490 20924 9496 20936
rect 9355 20896 9496 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 11609 20927 11667 20933
rect 11609 20924 11621 20927
rect 9600 20896 11621 20924
rect 4154 20856 4160 20868
rect 3252 20828 3832 20856
rect 3896 20828 4160 20856
rect 474 20748 480 20800
rect 532 20788 538 20800
rect 3252 20788 3280 20828
rect 532 20760 3280 20788
rect 532 20748 538 20760
rect 3602 20748 3608 20800
rect 3660 20748 3666 20800
rect 3804 20788 3832 20828
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 5644 20828 6500 20856
rect 5644 20788 5672 20828
rect 3804 20760 5672 20788
rect 5902 20748 5908 20800
rect 5960 20748 5966 20800
rect 6472 20788 6500 20828
rect 6546 20816 6552 20868
rect 6604 20816 6610 20868
rect 7558 20816 7564 20868
rect 7616 20816 7622 20868
rect 9600 20856 9628 20896
rect 11609 20893 11621 20896
rect 11655 20893 11667 20927
rect 11609 20887 11667 20893
rect 12161 20927 12219 20933
rect 12161 20893 12173 20927
rect 12207 20924 12219 20927
rect 12342 20924 12348 20936
rect 12207 20896 12348 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 7944 20828 9628 20856
rect 7944 20788 7972 20828
rect 9674 20816 9680 20868
rect 9732 20856 9738 20868
rect 10045 20859 10103 20865
rect 10045 20856 10057 20859
rect 9732 20828 10057 20856
rect 9732 20816 9738 20828
rect 10045 20825 10057 20828
rect 10091 20825 10103 20859
rect 10045 20819 10103 20825
rect 11057 20859 11115 20865
rect 11057 20825 11069 20859
rect 11103 20856 11115 20859
rect 11624 20856 11652 20887
rect 12342 20884 12348 20896
rect 12400 20924 12406 20936
rect 12636 20924 12664 20964
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 13817 20995 13875 21001
rect 13817 20961 13829 20995
rect 13863 20992 13875 20995
rect 14090 20992 14096 21004
rect 13863 20964 14096 20992
rect 13863 20961 13875 20964
rect 13817 20955 13875 20961
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 12400 20896 12664 20924
rect 12400 20884 12406 20896
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 14200 20924 14228 21032
rect 14274 20952 14280 21004
rect 14332 20952 14338 21004
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20992 14519 20995
rect 14918 20992 14924 21004
rect 14507 20964 14924 20992
rect 14507 20961 14519 20964
rect 14461 20955 14519 20961
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 15396 21001 15424 21032
rect 16408 21032 17408 21060
rect 15197 20995 15255 21001
rect 15197 20992 15209 20995
rect 15068 20964 15209 20992
rect 15068 20952 15074 20964
rect 15197 20961 15209 20964
rect 15243 20961 15255 20995
rect 15197 20955 15255 20961
rect 15381 20995 15439 21001
rect 15381 20961 15393 20995
rect 15427 20992 15439 20995
rect 15654 20992 15660 21004
rect 15427 20964 15660 20992
rect 15427 20961 15439 20964
rect 15381 20955 15439 20961
rect 15654 20952 15660 20964
rect 15712 20952 15718 21004
rect 16408 21001 16436 21032
rect 17402 21020 17408 21032
rect 17460 21020 17466 21072
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20961 16451 20995
rect 16393 20955 16451 20961
rect 16482 20952 16488 21004
rect 16540 20952 16546 21004
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17589 20995 17647 21001
rect 17589 20992 17601 20995
rect 17092 20964 17601 20992
rect 17092 20952 17098 20964
rect 17589 20961 17601 20964
rect 17635 20961 17647 20995
rect 17696 20992 17724 21100
rect 19061 21097 19073 21131
rect 19107 21128 19119 21131
rect 21818 21128 21824 21140
rect 19107 21100 21824 21128
rect 19107 21097 19119 21100
rect 19061 21091 19119 21097
rect 21818 21088 21824 21100
rect 21876 21088 21882 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 23017 21131 23075 21137
rect 23017 21128 23029 21131
rect 22336 21100 23029 21128
rect 22336 21088 22342 21100
rect 23017 21097 23029 21100
rect 23063 21097 23075 21131
rect 23017 21091 23075 21097
rect 25240 21100 27292 21128
rect 20714 21020 20720 21072
rect 20772 21060 20778 21072
rect 20772 21032 23704 21060
rect 20772 21020 20778 21032
rect 23676 21004 23704 21032
rect 19334 20992 19340 21004
rect 17696 20964 19340 20992
rect 17589 20955 17647 20961
rect 19334 20952 19340 20964
rect 19392 20952 19398 21004
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 20162 20992 20168 21004
rect 19484 20964 20168 20992
rect 19484 20952 19490 20964
rect 20162 20952 20168 20964
rect 20220 20992 20226 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 20220 20964 22385 20992
rect 20220 20952 20226 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 22462 20952 22468 21004
rect 22520 20992 22526 21004
rect 23477 20995 23535 21001
rect 23477 20992 23489 20995
rect 22520 20964 23489 20992
rect 22520 20952 22526 20964
rect 23477 20961 23489 20964
rect 23523 20961 23535 20995
rect 23477 20955 23535 20961
rect 23658 20952 23664 21004
rect 23716 20952 23722 21004
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20992 25191 20995
rect 25240 20992 25268 21100
rect 25958 21060 25964 21072
rect 25332 21032 25964 21060
rect 25332 21001 25360 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 27264 21060 27292 21100
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 27709 21131 27767 21137
rect 27709 21128 27721 21131
rect 27580 21100 27721 21128
rect 27580 21088 27586 21100
rect 27709 21097 27721 21100
rect 27755 21097 27767 21131
rect 27709 21091 27767 21097
rect 28902 21088 28908 21140
rect 28960 21128 28966 21140
rect 29273 21131 29331 21137
rect 29273 21128 29285 21131
rect 28960 21100 29285 21128
rect 28960 21088 28966 21100
rect 29273 21097 29285 21100
rect 29319 21097 29331 21131
rect 29273 21091 29331 21097
rect 31754 21088 31760 21140
rect 31812 21128 31818 21140
rect 31849 21131 31907 21137
rect 31849 21128 31861 21131
rect 31812 21100 31861 21128
rect 31812 21088 31818 21100
rect 31849 21097 31861 21100
rect 31895 21128 31907 21131
rect 32030 21128 32036 21140
rect 31895 21100 32036 21128
rect 31895 21097 31907 21100
rect 31849 21091 31907 21097
rect 32030 21088 32036 21100
rect 32088 21088 32094 21140
rect 33962 21088 33968 21140
rect 34020 21128 34026 21140
rect 34149 21131 34207 21137
rect 34149 21128 34161 21131
rect 34020 21100 34161 21128
rect 34020 21088 34026 21100
rect 34149 21097 34161 21100
rect 34195 21097 34207 21131
rect 34149 21091 34207 21097
rect 37366 21088 37372 21140
rect 37424 21088 37430 21140
rect 30650 21060 30656 21072
rect 27264 21032 30656 21060
rect 30650 21020 30656 21032
rect 30708 21020 30714 21072
rect 32398 21020 32404 21072
rect 32456 21060 32462 21072
rect 35897 21063 35955 21069
rect 35897 21060 35909 21063
rect 32456 21032 35909 21060
rect 32456 21020 32462 21032
rect 35897 21029 35909 21032
rect 35943 21029 35955 21063
rect 35897 21023 35955 21029
rect 25179 20964 25268 20992
rect 25317 20995 25375 21001
rect 25179 20961 25191 20964
rect 25133 20955 25191 20961
rect 25317 20961 25329 20995
rect 25363 20961 25375 20995
rect 26694 20992 26700 21004
rect 25317 20955 25375 20961
rect 25976 20964 26700 20992
rect 12768 20896 14228 20924
rect 12768 20884 12774 20896
rect 14826 20884 14832 20936
rect 14884 20924 14890 20936
rect 15105 20927 15163 20933
rect 15105 20924 15117 20927
rect 14884 20896 15117 20924
rect 14884 20884 14890 20896
rect 15105 20893 15117 20896
rect 15151 20893 15163 20927
rect 15105 20887 15163 20893
rect 16298 20884 16304 20936
rect 16356 20884 16362 20936
rect 17129 20927 17187 20933
rect 17129 20893 17141 20927
rect 17175 20893 17187 20927
rect 17129 20887 17187 20893
rect 17144 20856 17172 20887
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 19242 20924 19248 20936
rect 18564 20896 19248 20924
rect 18564 20884 18570 20896
rect 19242 20884 19248 20896
rect 19300 20884 19306 20936
rect 24302 20884 24308 20936
rect 24360 20924 24366 20936
rect 25976 20933 26004 20964
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 26970 20952 26976 21004
rect 27028 20992 27034 21004
rect 32217 20995 32275 21001
rect 32217 20992 32229 20995
rect 27028 20964 29776 20992
rect 27028 20952 27034 20964
rect 25961 20927 26019 20933
rect 25961 20924 25973 20927
rect 24360 20896 25973 20924
rect 24360 20884 24366 20896
rect 25961 20893 25973 20896
rect 26007 20893 26019 20927
rect 25961 20887 26019 20893
rect 28169 20927 28227 20933
rect 28169 20893 28181 20927
rect 28215 20924 28227 20927
rect 28442 20924 28448 20936
rect 28215 20896 28448 20924
rect 28215 20893 28227 20896
rect 28169 20887 28227 20893
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28534 20884 28540 20936
rect 28592 20924 28598 20936
rect 29086 20924 29092 20936
rect 28592 20896 29092 20924
rect 28592 20884 28598 20896
rect 29086 20884 29092 20896
rect 29144 20884 29150 20936
rect 29181 20927 29239 20933
rect 29181 20893 29193 20927
rect 29227 20924 29239 20927
rect 29362 20924 29368 20936
rect 29227 20896 29368 20924
rect 29227 20893 29239 20896
rect 29181 20887 29239 20893
rect 29362 20884 29368 20896
rect 29420 20884 29426 20936
rect 29748 20933 29776 20964
rect 31726 20964 32229 20992
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20924 29791 20927
rect 30190 20924 30196 20936
rect 29779 20896 30196 20924
rect 29779 20893 29791 20896
rect 29733 20887 29791 20893
rect 30190 20884 30196 20896
rect 30248 20884 30254 20936
rect 30834 20884 30840 20936
rect 30892 20884 30898 20936
rect 11103 20828 11560 20856
rect 11624 20828 17172 20856
rect 11103 20825 11115 20828
rect 11057 20819 11115 20825
rect 6472 20760 7972 20788
rect 8386 20748 8392 20800
rect 8444 20788 8450 20800
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 8444 20760 8493 20788
rect 8444 20748 8450 20760
rect 8481 20757 8493 20760
rect 8527 20788 8539 20791
rect 8570 20788 8576 20800
rect 8527 20760 8576 20788
rect 8527 20757 8539 20760
rect 8481 20751 8539 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 11146 20748 11152 20800
rect 11204 20748 11210 20800
rect 11532 20788 11560 20828
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 19260 20856 19288 20884
rect 19610 20856 19616 20868
rect 17276 20828 18920 20856
rect 19260 20828 19616 20856
rect 17276 20816 17282 20828
rect 12250 20788 12256 20800
rect 11532 20760 12256 20788
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 13906 20788 13912 20800
rect 12400 20760 13912 20788
rect 12400 20748 12406 20760
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14734 20748 14740 20800
rect 14792 20748 14798 20800
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16390 20788 16396 20800
rect 15979 20760 16396 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16390 20748 16396 20760
rect 16448 20748 16454 20800
rect 18782 20748 18788 20800
rect 18840 20748 18846 20800
rect 18892 20788 18920 20828
rect 19610 20816 19616 20828
rect 19668 20816 19674 20868
rect 19712 20859 19770 20865
rect 19712 20825 19724 20859
rect 19758 20856 19770 20859
rect 19758 20828 19932 20856
rect 19758 20825 19770 20828
rect 19712 20819 19770 20825
rect 19426 20788 19432 20800
rect 18892 20760 19432 20788
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 19904 20788 19932 20828
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 20036 20828 20194 20856
rect 20036 20816 20042 20828
rect 21634 20816 21640 20868
rect 21692 20816 21698 20868
rect 21818 20816 21824 20868
rect 21876 20856 21882 20868
rect 23385 20859 23443 20865
rect 23385 20856 23397 20859
rect 21876 20828 23397 20856
rect 21876 20816 21882 20828
rect 23385 20825 23397 20828
rect 23431 20856 23443 20859
rect 23750 20856 23756 20868
rect 23431 20828 23756 20856
rect 23431 20825 23443 20828
rect 23385 20819 23443 20825
rect 23750 20816 23756 20828
rect 23808 20816 23814 20868
rect 23934 20816 23940 20868
rect 23992 20856 23998 20868
rect 24854 20856 24860 20868
rect 23992 20828 24860 20856
rect 23992 20816 23998 20828
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 25087 20828 26188 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 20346 20788 20352 20800
rect 19904 20760 20352 20788
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 21082 20748 21088 20800
rect 21140 20788 21146 20800
rect 21177 20791 21235 20797
rect 21177 20788 21189 20791
rect 21140 20760 21189 20788
rect 21140 20748 21146 20760
rect 21177 20757 21189 20760
rect 21223 20757 21235 20791
rect 21177 20751 21235 20757
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 24213 20791 24271 20797
rect 24213 20788 24225 20791
rect 23624 20760 24225 20788
rect 23624 20748 23630 20760
rect 24213 20757 24225 20760
rect 24259 20788 24271 20791
rect 24302 20788 24308 20800
rect 24259 20760 24308 20788
rect 24259 20757 24271 20760
rect 24213 20751 24271 20757
rect 24302 20748 24308 20760
rect 24360 20748 24366 20800
rect 24578 20748 24584 20800
rect 24636 20788 24642 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 24636 20760 24685 20788
rect 24636 20748 24642 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24872 20788 24900 20816
rect 25590 20788 25596 20800
rect 24872 20760 25596 20788
rect 24673 20751 24731 20757
rect 25590 20748 25596 20760
rect 25648 20748 25654 20800
rect 26160 20788 26188 20828
rect 26234 20816 26240 20868
rect 26292 20816 26298 20868
rect 26510 20816 26516 20868
rect 26568 20856 26574 20868
rect 31726 20856 31754 20964
rect 32217 20961 32229 20964
rect 32263 20961 32275 20995
rect 32217 20955 32275 20961
rect 32858 20952 32864 21004
rect 32916 20952 32922 21004
rect 33137 20995 33195 21001
rect 33137 20961 33149 20995
rect 33183 20992 33195 20995
rect 33318 20992 33324 21004
rect 33183 20964 33324 20992
rect 33183 20961 33195 20964
rect 33137 20955 33195 20961
rect 33318 20952 33324 20964
rect 33376 20952 33382 21004
rect 34330 20884 34336 20936
rect 34388 20884 34394 20936
rect 36630 20884 36636 20936
rect 36688 20924 36694 20936
rect 46842 20924 46848 20936
rect 36688 20896 46848 20924
rect 36688 20884 36694 20896
rect 46842 20884 46848 20896
rect 46900 20884 46906 20936
rect 26568 20828 26726 20856
rect 27632 20828 31754 20856
rect 34977 20859 35035 20865
rect 26568 20816 26574 20828
rect 27632 20788 27660 20828
rect 34977 20825 34989 20859
rect 35023 20856 35035 20859
rect 35250 20856 35256 20868
rect 35023 20828 35256 20856
rect 35023 20825 35035 20828
rect 34977 20819 35035 20825
rect 35250 20816 35256 20828
rect 35308 20816 35314 20868
rect 35434 20816 35440 20868
rect 35492 20856 35498 20868
rect 35713 20859 35771 20865
rect 35713 20856 35725 20859
rect 35492 20828 35725 20856
rect 35492 20816 35498 20828
rect 35713 20825 35725 20828
rect 35759 20825 35771 20859
rect 35713 20819 35771 20825
rect 36446 20816 36452 20868
rect 36504 20856 36510 20868
rect 36909 20859 36967 20865
rect 36909 20856 36921 20859
rect 36504 20828 36921 20856
rect 36504 20816 36510 20828
rect 36909 20825 36921 20828
rect 36955 20825 36967 20859
rect 36909 20819 36967 20825
rect 26160 20760 27660 20788
rect 28810 20748 28816 20800
rect 28868 20748 28874 20800
rect 29178 20748 29184 20800
rect 29236 20788 29242 20800
rect 30377 20791 30435 20797
rect 30377 20788 30389 20791
rect 29236 20760 30389 20788
rect 29236 20748 29242 20760
rect 30377 20757 30389 20760
rect 30423 20757 30435 20791
rect 30377 20751 30435 20757
rect 31478 20748 31484 20800
rect 31536 20748 31542 20800
rect 35066 20748 35072 20800
rect 35124 20748 35130 20800
rect 36538 20748 36544 20800
rect 36596 20748 36602 20800
rect 37090 20748 37096 20800
rect 37148 20748 37154 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 1026 20544 1032 20596
rect 1084 20584 1090 20596
rect 5258 20584 5264 20596
rect 1084 20556 5264 20584
rect 1084 20544 1090 20556
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 6454 20584 6460 20596
rect 5675 20556 6460 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 11057 20587 11115 20593
rect 11057 20584 11069 20587
rect 7116 20556 11069 20584
rect 6178 20516 6184 20528
rect 3620 20488 6184 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 1946 20448 1952 20460
rect 1811 20420 1952 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 3620 20457 3648 20488
rect 6178 20476 6184 20488
rect 6236 20476 6242 20528
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 5626 20448 5632 20460
rect 3605 20411 3663 20417
rect 3804 20420 5632 20448
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3804 20380 3832 20420
rect 5626 20408 5632 20420
rect 5684 20408 5690 20460
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20448 5779 20451
rect 6362 20448 6368 20460
rect 5767 20420 6368 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 3620 20352 3832 20380
rect 2406 20272 2412 20324
rect 2464 20312 2470 20324
rect 3620 20312 3648 20352
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5813 20383 5871 20389
rect 5813 20380 5825 20383
rect 5592 20352 5825 20380
rect 5592 20340 5598 20352
rect 5813 20349 5825 20352
rect 5859 20349 5871 20383
rect 5813 20343 5871 20349
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 6564 20380 6592 20411
rect 5960 20352 6592 20380
rect 5960 20340 5966 20352
rect 6638 20340 6644 20392
rect 6696 20380 6702 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 6696 20352 7021 20380
rect 6696 20340 6702 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 2464 20284 3648 20312
rect 2464 20272 2470 20284
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 7116 20312 7144 20556
rect 11057 20553 11069 20556
rect 11103 20553 11115 20587
rect 11057 20547 11115 20553
rect 11974 20544 11980 20596
rect 12032 20544 12038 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 15562 20584 15568 20596
rect 13035 20556 15568 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 16942 20584 16948 20596
rect 16724 20556 16948 20584
rect 16724 20544 16730 20556
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17494 20544 17500 20596
rect 17552 20544 17558 20596
rect 18141 20587 18199 20593
rect 18141 20584 18153 20587
rect 17696 20556 18153 20584
rect 9122 20516 9128 20528
rect 8312 20488 9128 20516
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 8312 20389 8340 20488
rect 9122 20476 9128 20488
rect 9180 20516 9186 20528
rect 9180 20488 9338 20516
rect 9180 20476 9186 20488
rect 11238 20476 11244 20528
rect 11296 20516 11302 20528
rect 11698 20516 11704 20528
rect 11296 20488 11704 20516
rect 11296 20476 11302 20488
rect 11698 20476 11704 20488
rect 11756 20516 11762 20528
rect 11885 20519 11943 20525
rect 11885 20516 11897 20519
rect 11756 20488 11897 20516
rect 11756 20476 11762 20488
rect 11885 20485 11897 20488
rect 11931 20485 11943 20519
rect 11885 20479 11943 20485
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 12897 20519 12955 20525
rect 12897 20516 12909 20519
rect 12860 20488 12909 20516
rect 12860 20476 12866 20488
rect 12897 20485 12909 20488
rect 12943 20516 12955 20519
rect 13630 20516 13636 20528
rect 12943 20488 13636 20516
rect 12943 20485 12955 20488
rect 12897 20479 12955 20485
rect 13630 20476 13636 20488
rect 13688 20476 13694 20528
rect 13998 20476 14004 20528
rect 14056 20516 14062 20528
rect 14274 20516 14280 20528
rect 14056 20488 14280 20516
rect 14056 20476 14062 20488
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 14550 20476 14556 20528
rect 14608 20476 14614 20528
rect 16960 20516 16988 20544
rect 17696 20516 17724 20556
rect 18141 20553 18153 20556
rect 18187 20553 18199 20587
rect 18141 20547 18199 20553
rect 18966 20544 18972 20596
rect 19024 20544 19030 20596
rect 20364 20556 21312 20584
rect 16960 20488 17724 20516
rect 17770 20476 17776 20528
rect 17828 20516 17834 20528
rect 20364 20516 20392 20556
rect 17828 20488 20392 20516
rect 17828 20476 17834 20488
rect 20714 20476 20720 20528
rect 20772 20476 20778 20528
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10744 20420 10977 20448
rect 10744 20408 10750 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 13538 20448 13544 20460
rect 10965 20411 11023 20417
rect 13004 20420 13544 20448
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 7616 20352 8309 20380
rect 7616 20340 7622 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 8573 20383 8631 20389
rect 8573 20349 8585 20383
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 3752 20284 7144 20312
rect 3752 20272 3758 20284
rect 7282 20272 7288 20324
rect 7340 20312 7346 20324
rect 7834 20312 7840 20324
rect 7340 20284 7840 20312
rect 7340 20272 7346 20284
rect 7834 20272 7840 20284
rect 7892 20312 7898 20324
rect 8588 20312 8616 20343
rect 8846 20340 8852 20392
rect 8904 20340 8910 20392
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 10321 20383 10379 20389
rect 10321 20380 10333 20383
rect 9548 20352 10333 20380
rect 9548 20340 9554 20352
rect 10321 20349 10333 20352
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 13004 20380 13032 20420
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13722 20408 13728 20460
rect 13780 20408 13786 20460
rect 16022 20408 16028 20460
rect 16080 20408 16086 20460
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20448 17463 20451
rect 17862 20448 17868 20460
rect 17451 20420 17868 20448
rect 17451 20417 17463 20420
rect 17405 20411 17463 20417
rect 17862 20408 17868 20420
rect 17920 20408 17926 20460
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 18877 20451 18935 20457
rect 18877 20448 18889 20451
rect 18840 20420 18889 20448
rect 18840 20408 18846 20420
rect 18877 20417 18889 20420
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 18984 20420 19288 20448
rect 10928 20352 13032 20380
rect 13173 20383 13231 20389
rect 10928 20340 10934 20352
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13354 20380 13360 20392
rect 13219 20352 13360 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13354 20340 13360 20352
rect 13412 20340 13418 20392
rect 14090 20340 14096 20392
rect 14148 20380 14154 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 14148 20352 15485 20380
rect 14148 20340 14154 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 17589 20383 17647 20389
rect 17589 20380 17601 20383
rect 15473 20343 15531 20349
rect 16960 20352 17601 20380
rect 7892 20284 8616 20312
rect 7892 20272 7898 20284
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 5718 20244 5724 20256
rect 5307 20216 5724 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 5810 20204 5816 20256
rect 5868 20244 5874 20256
rect 8202 20244 8208 20256
rect 5868 20216 8208 20244
rect 5868 20204 5874 20216
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8588 20244 8616 20284
rect 9950 20272 9956 20324
rect 10008 20312 10014 20324
rect 16209 20315 16267 20321
rect 16209 20312 16221 20315
rect 10008 20284 13860 20312
rect 10008 20272 10014 20284
rect 9398 20244 9404 20256
rect 8588 20216 9404 20244
rect 9398 20204 9404 20216
rect 9456 20244 9462 20256
rect 9858 20244 9864 20256
rect 9456 20216 9864 20244
rect 9456 20204 9462 20216
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11422 20244 11428 20256
rect 11112 20216 11428 20244
rect 11112 20204 11118 20216
rect 11422 20204 11428 20216
rect 11480 20244 11486 20256
rect 12342 20244 12348 20256
rect 11480 20216 12348 20244
rect 11480 20204 11486 20216
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 12529 20247 12587 20253
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 12710 20244 12716 20256
rect 12575 20216 12716 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13832 20244 13860 20284
rect 15028 20284 16221 20312
rect 15028 20244 15056 20284
rect 16209 20281 16221 20284
rect 16255 20281 16267 20315
rect 16209 20275 16267 20281
rect 13832 20216 15056 20244
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 16960 20244 16988 20352
rect 17589 20349 17601 20352
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 17604 20312 17632 20343
rect 17678 20340 17684 20392
rect 17736 20380 17742 20392
rect 18984 20380 19012 20420
rect 17736 20352 19012 20380
rect 17736 20340 17742 20352
rect 19150 20340 19156 20392
rect 19208 20340 19214 20392
rect 19260 20380 19288 20420
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19668 20420 19717 20448
rect 19668 20408 19674 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 21284 20448 21312 20556
rect 23566 20544 23572 20596
rect 23624 20544 23630 20596
rect 23842 20544 23848 20596
rect 23900 20584 23906 20596
rect 27157 20587 27215 20593
rect 27157 20584 27169 20587
rect 23900 20556 27169 20584
rect 23900 20544 23906 20556
rect 27157 20553 27169 20556
rect 27203 20553 27215 20587
rect 27157 20547 27215 20553
rect 27430 20544 27436 20596
rect 27488 20584 27494 20596
rect 31478 20584 31484 20596
rect 27488 20556 27844 20584
rect 27488 20544 27494 20556
rect 23382 20476 23388 20528
rect 23440 20516 23446 20528
rect 23477 20519 23535 20525
rect 23477 20516 23489 20519
rect 23440 20488 23489 20516
rect 23440 20476 23446 20488
rect 23477 20485 23489 20488
rect 23523 20516 23535 20519
rect 23523 20488 24256 20516
rect 23523 20485 23535 20488
rect 23477 20479 23535 20485
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21284 20420 22017 20448
rect 19705 20411 19763 20417
rect 22005 20417 22017 20420
rect 22051 20448 22063 20451
rect 22051 20420 23520 20448
rect 22051 20417 22063 20420
rect 22005 20411 22063 20417
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 19260 20352 21465 20380
rect 21453 20349 21465 20352
rect 21499 20380 21511 20383
rect 23382 20380 23388 20392
rect 21499 20352 23388 20380
rect 21499 20349 21511 20352
rect 21453 20343 21511 20349
rect 23382 20340 23388 20352
rect 23440 20340 23446 20392
rect 19702 20312 19708 20324
rect 17604 20284 19708 20312
rect 19702 20272 19708 20284
rect 19760 20272 19766 20324
rect 20990 20272 20996 20324
rect 21048 20312 21054 20324
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 21048 20284 23121 20312
rect 21048 20272 21054 20284
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 15252 20216 16988 20244
rect 15252 20204 15258 20216
rect 17034 20204 17040 20256
rect 17092 20204 17098 20256
rect 17126 20204 17132 20256
rect 17184 20244 17190 20256
rect 18230 20244 18236 20256
rect 17184 20216 18236 20244
rect 17184 20204 17190 20216
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 18414 20204 18420 20256
rect 18472 20244 18478 20256
rect 18509 20247 18567 20253
rect 18509 20244 18521 20247
rect 18472 20216 18521 20244
rect 18472 20204 18478 20216
rect 18509 20213 18521 20216
rect 18555 20213 18567 20247
rect 18509 20207 18567 20213
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 19962 20247 20020 20253
rect 19962 20244 19974 20247
rect 18748 20216 19974 20244
rect 18748 20204 18754 20216
rect 19962 20213 19974 20216
rect 20008 20213 20020 20247
rect 19962 20207 20020 20213
rect 22646 20204 22652 20256
rect 22704 20204 22710 20256
rect 23492 20244 23520 20420
rect 23750 20340 23756 20392
rect 23808 20340 23814 20392
rect 24228 20312 24256 20488
rect 24486 20476 24492 20528
rect 24544 20516 24550 20528
rect 24581 20519 24639 20525
rect 24581 20516 24593 20519
rect 24544 20488 24593 20516
rect 24544 20476 24550 20488
rect 24581 20485 24593 20488
rect 24627 20485 24639 20519
rect 24581 20479 24639 20485
rect 24854 20476 24860 20528
rect 24912 20516 24918 20528
rect 26421 20519 26479 20525
rect 24912 20488 25070 20516
rect 24912 20476 24918 20488
rect 26421 20485 26433 20519
rect 26467 20516 26479 20519
rect 26510 20516 26516 20528
rect 26467 20488 26516 20516
rect 26467 20485 26479 20488
rect 26421 20479 26479 20485
rect 26510 20476 26516 20488
rect 26568 20516 26574 20528
rect 26878 20516 26884 20528
rect 26568 20488 26884 20516
rect 26568 20476 26574 20488
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 26970 20476 26976 20528
rect 27028 20516 27034 20528
rect 27028 20488 27752 20516
rect 27028 20476 27034 20488
rect 26789 20451 26847 20457
rect 26789 20417 26801 20451
rect 26835 20448 26847 20451
rect 27522 20448 27528 20460
rect 26835 20420 27528 20448
rect 26835 20417 26847 20420
rect 26789 20411 26847 20417
rect 24302 20340 24308 20392
rect 24360 20340 24366 20392
rect 25314 20380 25320 20392
rect 24412 20352 25320 20380
rect 24412 20312 24440 20352
rect 25314 20340 25320 20352
rect 25372 20380 25378 20392
rect 26804 20380 26832 20411
rect 27522 20408 27528 20420
rect 27580 20408 27586 20460
rect 25372 20352 26832 20380
rect 25372 20340 25378 20352
rect 27154 20340 27160 20392
rect 27212 20380 27218 20392
rect 27724 20389 27752 20488
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 27212 20352 27629 20380
rect 27212 20340 27218 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27709 20383 27767 20389
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27816 20380 27844 20556
rect 28736 20556 31484 20584
rect 28736 20525 28764 20556
rect 31478 20544 31484 20556
rect 31536 20544 31542 20596
rect 31754 20544 31760 20596
rect 31812 20544 31818 20596
rect 31846 20544 31852 20596
rect 31904 20544 31910 20596
rect 32858 20544 32864 20596
rect 32916 20584 32922 20596
rect 33229 20587 33287 20593
rect 33229 20584 33241 20587
rect 32916 20556 33241 20584
rect 32916 20544 32922 20556
rect 33229 20553 33241 20556
rect 33275 20553 33287 20587
rect 33229 20547 33287 20553
rect 34974 20544 34980 20596
rect 35032 20584 35038 20596
rect 35032 20556 35204 20584
rect 35032 20544 35038 20556
rect 28721 20519 28779 20525
rect 28721 20485 28733 20519
rect 28767 20485 28779 20519
rect 28721 20479 28779 20485
rect 29362 20476 29368 20528
rect 29420 20476 29426 20528
rect 30024 20488 32628 20516
rect 27982 20408 27988 20460
rect 28040 20448 28046 20460
rect 28350 20448 28356 20460
rect 28040 20420 28356 20448
rect 28040 20408 28046 20420
rect 28350 20408 28356 20420
rect 28408 20448 28414 20460
rect 28445 20451 28503 20457
rect 28445 20448 28457 20451
rect 28408 20420 28457 20448
rect 28408 20408 28414 20420
rect 28445 20417 28457 20420
rect 28491 20417 28503 20451
rect 28445 20411 28503 20417
rect 30024 20380 30052 20488
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 31113 20451 31171 20457
rect 31113 20417 31125 20451
rect 31159 20448 31171 20451
rect 31159 20420 32260 20448
rect 31159 20417 31171 20420
rect 31113 20411 31171 20417
rect 27816 20352 30052 20380
rect 27709 20343 27767 20349
rect 24228 20284 24440 20312
rect 26053 20315 26111 20321
rect 26053 20281 26065 20315
rect 26099 20312 26111 20315
rect 26970 20312 26976 20324
rect 26099 20284 26976 20312
rect 26099 20281 26111 20284
rect 26053 20275 26111 20281
rect 26970 20272 26976 20284
rect 27028 20272 27034 20324
rect 27724 20312 27752 20343
rect 30190 20340 30196 20392
rect 30248 20340 30254 20392
rect 28074 20312 28080 20324
rect 27724 20284 28080 20312
rect 28074 20272 28080 20284
rect 28132 20272 28138 20324
rect 30374 20312 30380 20324
rect 29840 20284 30380 20312
rect 24762 20244 24768 20256
rect 23492 20216 24768 20244
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 26513 20247 26571 20253
rect 26513 20244 26525 20247
rect 26292 20216 26525 20244
rect 26292 20204 26298 20216
rect 26513 20213 26525 20216
rect 26559 20213 26571 20247
rect 26513 20207 26571 20213
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 29840 20244 29868 20284
rect 30374 20272 30380 20284
rect 30432 20272 30438 20324
rect 31036 20312 31064 20411
rect 31202 20340 31208 20392
rect 31260 20340 31266 20392
rect 31846 20312 31852 20324
rect 31036 20284 31852 20312
rect 31846 20272 31852 20284
rect 31904 20272 31910 20324
rect 32232 20312 32260 20420
rect 32306 20408 32312 20460
rect 32364 20408 32370 20460
rect 32600 20380 32628 20488
rect 32674 20476 32680 20528
rect 32732 20516 32738 20528
rect 34425 20519 34483 20525
rect 34425 20516 34437 20519
rect 32732 20488 34437 20516
rect 32732 20476 32738 20488
rect 34425 20485 34437 20488
rect 34471 20516 34483 20519
rect 35069 20519 35127 20525
rect 35069 20516 35081 20519
rect 34471 20488 35081 20516
rect 34471 20485 34483 20488
rect 34425 20479 34483 20485
rect 35069 20485 35081 20488
rect 35115 20485 35127 20519
rect 35176 20516 35204 20556
rect 35526 20544 35532 20596
rect 35584 20584 35590 20596
rect 35621 20587 35679 20593
rect 35621 20584 35633 20587
rect 35584 20556 35633 20584
rect 35584 20544 35590 20556
rect 35621 20553 35633 20556
rect 35667 20553 35679 20587
rect 35621 20547 35679 20553
rect 39574 20516 39580 20528
rect 35176 20488 39580 20516
rect 35069 20479 35127 20485
rect 39574 20476 39580 20488
rect 39632 20476 39638 20528
rect 33686 20408 33692 20460
rect 33744 20448 33750 20460
rect 34885 20451 34943 20457
rect 34885 20448 34897 20451
rect 33744 20420 34897 20448
rect 33744 20408 33750 20420
rect 34885 20417 34897 20420
rect 34931 20417 34943 20451
rect 40954 20448 40960 20460
rect 34885 20411 34943 20417
rect 34992 20420 40960 20448
rect 34992 20380 35020 20420
rect 40954 20408 40960 20420
rect 41012 20408 41018 20460
rect 35618 20380 35624 20392
rect 32600 20352 35020 20380
rect 35268 20352 35624 20380
rect 34974 20312 34980 20324
rect 32232 20284 34980 20312
rect 34974 20272 34980 20284
rect 35032 20272 35038 20324
rect 35158 20272 35164 20324
rect 35216 20312 35222 20324
rect 35268 20312 35296 20352
rect 35618 20340 35624 20352
rect 35676 20380 35682 20392
rect 35989 20383 36047 20389
rect 35989 20380 36001 20383
rect 35676 20352 36001 20380
rect 35676 20340 35682 20352
rect 35989 20349 36001 20352
rect 36035 20349 36047 20383
rect 35989 20343 36047 20349
rect 35216 20284 35296 20312
rect 35216 20272 35222 20284
rect 35342 20272 35348 20324
rect 35400 20312 35406 20324
rect 35710 20312 35716 20324
rect 35400 20284 35716 20312
rect 35400 20272 35406 20284
rect 35710 20272 35716 20284
rect 35768 20312 35774 20324
rect 35897 20315 35955 20321
rect 35897 20312 35909 20315
rect 35768 20284 35909 20312
rect 35768 20272 35774 20284
rect 35897 20281 35909 20284
rect 35943 20281 35955 20315
rect 35897 20275 35955 20281
rect 27580 20216 29868 20244
rect 27580 20204 27586 20216
rect 29914 20204 29920 20256
rect 29972 20244 29978 20256
rect 30653 20247 30711 20253
rect 30653 20244 30665 20247
rect 29972 20216 30665 20244
rect 29972 20204 29978 20216
rect 30653 20213 30665 20216
rect 30699 20213 30711 20247
rect 30653 20207 30711 20213
rect 32030 20204 32036 20256
rect 32088 20244 32094 20256
rect 32953 20247 33011 20253
rect 32953 20244 32965 20247
rect 32088 20216 32965 20244
rect 32088 20204 32094 20216
rect 32953 20213 32965 20216
rect 32999 20213 33011 20247
rect 32953 20207 33011 20213
rect 33778 20204 33784 20256
rect 33836 20204 33842 20256
rect 34514 20204 34520 20256
rect 34572 20204 34578 20256
rect 35250 20204 35256 20256
rect 35308 20204 35314 20256
rect 35434 20204 35440 20256
rect 35492 20204 35498 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3602 20000 3608 20052
rect 3660 20000 3666 20052
rect 4154 20000 4160 20052
rect 4212 20000 4218 20052
rect 6914 20040 6920 20052
rect 5000 20012 6920 20040
rect 3881 19975 3939 19981
rect 3881 19941 3893 19975
rect 3927 19972 3939 19975
rect 5000 19972 5028 20012
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 8941 20043 8999 20049
rect 8941 20040 8953 20043
rect 8260 20012 8953 20040
rect 8260 20000 8266 20012
rect 8941 20009 8953 20012
rect 8987 20040 8999 20043
rect 11606 20040 11612 20052
rect 8987 20012 11612 20040
rect 8987 20009 8999 20012
rect 8941 20003 8999 20009
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 14090 20040 14096 20052
rect 13372 20012 14096 20040
rect 3927 19944 5028 19972
rect 3927 19941 3939 19944
rect 3881 19935 3939 19941
rect 7834 19932 7840 19984
rect 7892 19972 7898 19984
rect 9490 19972 9496 19984
rect 7892 19944 9496 19972
rect 7892 19932 7898 19944
rect 9490 19932 9496 19944
rect 9548 19932 9554 19984
rect 11330 19932 11336 19984
rect 11388 19972 11394 19984
rect 13372 19972 13400 20012
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 15010 20040 15016 20052
rect 14608 20012 15016 20040
rect 14608 20000 14614 20012
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 15562 20000 15568 20052
rect 15620 20040 15626 20052
rect 15620 20012 16436 20040
rect 15620 20000 15626 20012
rect 13722 19972 13728 19984
rect 11388 19944 13400 19972
rect 13464 19944 13728 19972
rect 11388 19932 11394 19944
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 7374 19904 7380 19916
rect 3467 19876 7380 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 7374 19864 7380 19876
rect 7432 19864 7438 19916
rect 7466 19864 7472 19916
rect 7524 19904 7530 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 7524 19876 7573 19904
rect 7524 19864 7530 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 9950 19904 9956 19916
rect 7561 19867 7619 19873
rect 9324 19876 9956 19904
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19836 1823 19839
rect 2498 19836 2504 19848
rect 1811 19808 2504 19836
rect 1811 19805 1823 19808
rect 1765 19799 1823 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 2777 19771 2835 19777
rect 2777 19737 2789 19771
rect 2823 19768 2835 19771
rect 2866 19768 2872 19780
rect 2823 19740 2872 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 4356 19700 4384 19799
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 9324 19836 9352 19876
rect 9950 19864 9956 19876
rect 10008 19864 10014 19916
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19904 10103 19907
rect 13464 19904 13492 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 16408 19981 16436 20012
rect 17678 20000 17684 20052
rect 17736 20000 17742 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 18064 20012 18153 20040
rect 14185 19975 14243 19981
rect 14185 19941 14197 19975
rect 14231 19972 14243 19975
rect 16393 19975 16451 19981
rect 14231 19944 14780 19972
rect 14231 19941 14243 19944
rect 14185 19935 14243 19941
rect 10091 19876 13492 19904
rect 13633 19907 13691 19913
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 13633 19873 13645 19907
rect 13679 19873 13691 19907
rect 13740 19904 13768 19932
rect 14645 19907 14703 19913
rect 14645 19904 14657 19907
rect 13740 19876 14657 19904
rect 13633 19867 13691 19873
rect 14645 19873 14657 19876
rect 14691 19873 14703 19907
rect 14752 19904 14780 19944
rect 16393 19941 16405 19975
rect 16439 19972 16451 19975
rect 17126 19972 17132 19984
rect 16439 19944 17132 19972
rect 16439 19941 16451 19944
rect 16393 19935 16451 19941
rect 17126 19932 17132 19944
rect 17184 19932 17190 19984
rect 14752 19876 17724 19904
rect 14645 19867 14703 19873
rect 7331 19808 9352 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 9398 19796 9404 19848
rect 9456 19796 9462 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 13648 19836 13676 19867
rect 14090 19836 14096 19848
rect 11664 19808 13308 19836
rect 13648 19808 14096 19836
rect 11664 19796 11670 19808
rect 4522 19728 4528 19780
rect 4580 19768 4586 19780
rect 5169 19771 5227 19777
rect 5169 19768 5181 19771
rect 4580 19740 5181 19768
rect 4580 19728 4586 19740
rect 5169 19737 5181 19740
rect 5215 19737 5227 19771
rect 5169 19731 5227 19737
rect 5626 19728 5632 19780
rect 5684 19728 5690 19780
rect 8294 19728 8300 19780
rect 8352 19768 8358 19780
rect 8352 19740 9996 19768
rect 8352 19728 8358 19740
rect 5810 19700 5816 19712
rect 4356 19672 5816 19700
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6641 19703 6699 19709
rect 6641 19700 6653 19703
rect 6052 19672 6653 19700
rect 6052 19660 6058 19672
rect 6641 19669 6653 19672
rect 6687 19669 6699 19703
rect 6641 19663 6699 19669
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 6788 19672 9505 19700
rect 6788 19660 6794 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 9968 19700 9996 19740
rect 10042 19728 10048 19780
rect 10100 19768 10106 19780
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 10100 19740 10333 19768
rect 10100 19728 10106 19740
rect 10321 19737 10333 19740
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 11054 19728 11060 19780
rect 11112 19728 11118 19780
rect 12342 19728 12348 19780
rect 12400 19728 12406 19780
rect 12529 19771 12587 19777
rect 12529 19737 12541 19771
rect 12575 19768 12587 19771
rect 12802 19768 12808 19780
rect 12575 19740 12808 19768
rect 12575 19737 12587 19740
rect 12529 19731 12587 19737
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 13280 19768 13308 19808
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17126 19836 17132 19848
rect 17083 19808 17132 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17696 19836 17724 19876
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18064 19904 18092 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 20622 20040 20628 20052
rect 18141 20003 18199 20009
rect 19536 20012 20628 20040
rect 18230 19932 18236 19984
rect 18288 19972 18294 19984
rect 19426 19972 19432 19984
rect 18288 19944 19432 19972
rect 18288 19932 18294 19944
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18012 19876 18092 19904
rect 18248 19876 18705 19904
rect 18012 19864 18018 19876
rect 18248 19836 18276 19876
rect 18693 19873 18705 19876
rect 18739 19904 18751 19907
rect 19536 19904 19564 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21910 20000 21916 20052
rect 21968 20000 21974 20052
rect 22373 20043 22431 20049
rect 22373 20009 22385 20043
rect 22419 20040 22431 20043
rect 25958 20040 25964 20052
rect 22419 20012 25964 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 25958 20000 25964 20012
rect 26016 20000 26022 20052
rect 26132 20043 26190 20049
rect 26132 20009 26144 20043
rect 26178 20040 26190 20043
rect 27617 20043 27675 20049
rect 26178 20012 27476 20040
rect 26178 20009 26190 20012
rect 26132 20003 26190 20009
rect 27448 19972 27476 20012
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 27798 20040 27804 20052
rect 27663 20012 27804 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 27890 20000 27896 20052
rect 27948 20040 27954 20052
rect 27948 20012 31432 20040
rect 27948 20000 27954 20012
rect 28810 19972 28816 19984
rect 27448 19944 28816 19972
rect 28810 19932 28816 19944
rect 28868 19932 28874 19984
rect 28902 19932 28908 19984
rect 28960 19972 28966 19984
rect 31294 19972 31300 19984
rect 28960 19944 31300 19972
rect 28960 19932 28966 19944
rect 31294 19932 31300 19944
rect 31352 19932 31358 19984
rect 18739 19876 19564 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 19668 19876 19717 19904
rect 19668 19864 19674 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20441 19907 20499 19913
rect 20441 19873 20453 19907
rect 20487 19904 20499 19907
rect 22646 19904 22652 19916
rect 20487 19876 22652 19904
rect 20487 19873 20499 19876
rect 20441 19867 20499 19873
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 23661 19907 23719 19913
rect 23661 19873 23673 19907
rect 23707 19904 23719 19907
rect 25038 19904 25044 19916
rect 23707 19876 25044 19904
rect 23707 19873 23719 19876
rect 23661 19867 23719 19873
rect 25038 19864 25044 19876
rect 25096 19864 25102 19916
rect 25314 19864 25320 19916
rect 25372 19864 25378 19916
rect 25774 19864 25780 19916
rect 25832 19904 25838 19916
rect 25869 19907 25927 19913
rect 25869 19904 25881 19907
rect 25832 19876 25881 19904
rect 25832 19864 25838 19876
rect 25869 19873 25881 19876
rect 25915 19904 25927 19907
rect 27614 19904 27620 19916
rect 25915 19876 27620 19904
rect 25915 19873 25927 19876
rect 25869 19867 25927 19873
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 27706 19864 27712 19916
rect 27764 19904 27770 19916
rect 27764 19876 28212 19904
rect 27764 19864 27770 19876
rect 17696 19808 18276 19836
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 20070 19836 20076 19848
rect 18647 19808 20076 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 22554 19796 22560 19848
rect 22612 19796 22618 19848
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 23385 19839 23443 19845
rect 23385 19836 23397 19839
rect 22796 19808 23397 19836
rect 22796 19796 22802 19808
rect 23385 19805 23397 19808
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19836 23535 19839
rect 27632 19836 27660 19864
rect 27982 19836 27988 19848
rect 23523 19808 25360 19836
rect 27632 19808 27988 19836
rect 23523 19805 23535 19808
rect 23477 19799 23535 19805
rect 14921 19771 14979 19777
rect 14921 19768 14933 19771
rect 13280 19740 14933 19768
rect 14921 19737 14933 19740
rect 14967 19737 14979 19771
rect 14921 19731 14979 19737
rect 15010 19728 15016 19780
rect 15068 19768 15074 19780
rect 16666 19768 16672 19780
rect 15068 19740 15410 19768
rect 16408 19740 16672 19768
rect 15068 19728 15074 19740
rect 11330 19700 11336 19712
rect 9968 19672 11336 19700
rect 9493 19663 9551 19669
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 12250 19700 12256 19712
rect 11839 19672 12256 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 13354 19660 13360 19712
rect 13412 19660 13418 19712
rect 13446 19660 13452 19712
rect 13504 19660 13510 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 13998 19700 14004 19712
rect 13596 19672 14004 19700
rect 13596 19660 13602 19672
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 16408 19700 16436 19740
rect 16666 19728 16672 19740
rect 16724 19768 16730 19780
rect 18322 19768 18328 19780
rect 16724 19740 18328 19768
rect 16724 19728 16730 19740
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 18432 19740 19533 19768
rect 14415 19672 16436 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 16482 19660 16488 19712
rect 16540 19700 16546 19712
rect 18432 19700 18460 19740
rect 19521 19737 19533 19740
rect 19567 19768 19579 19771
rect 19886 19768 19892 19780
rect 19567 19740 19892 19768
rect 19567 19737 19579 19740
rect 19521 19731 19579 19737
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 20346 19728 20352 19780
rect 20404 19728 20410 19780
rect 20714 19728 20720 19780
rect 20772 19768 20778 19780
rect 25041 19771 25099 19777
rect 20772 19740 20930 19768
rect 22066 19740 24716 19768
rect 20772 19728 20778 19740
rect 16540 19672 18460 19700
rect 16540 19660 16546 19672
rect 18506 19660 18512 19712
rect 18564 19660 18570 19712
rect 19794 19660 19800 19712
rect 19852 19700 19858 19712
rect 20364 19700 20392 19728
rect 19852 19672 20392 19700
rect 19852 19660 19858 19672
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 22066 19700 22094 19740
rect 21140 19672 22094 19700
rect 21140 19660 21146 19672
rect 22922 19660 22928 19712
rect 22980 19700 22986 19712
rect 23017 19703 23075 19709
rect 23017 19700 23029 19703
rect 22980 19672 23029 19700
rect 22980 19660 22986 19672
rect 23017 19669 23029 19672
rect 23063 19669 23075 19703
rect 23017 19663 23075 19669
rect 23658 19660 23664 19712
rect 23716 19700 23722 19712
rect 24121 19703 24179 19709
rect 24121 19700 24133 19703
rect 23716 19672 24133 19700
rect 23716 19660 23722 19672
rect 24121 19669 24133 19672
rect 24167 19700 24179 19703
rect 24302 19700 24308 19712
rect 24167 19672 24308 19700
rect 24167 19669 24179 19672
rect 24121 19663 24179 19669
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 24688 19709 24716 19740
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 25222 19768 25228 19780
rect 25087 19740 25228 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 25332 19768 25360 19808
rect 27982 19796 27988 19808
rect 28040 19796 28046 19848
rect 28074 19796 28080 19848
rect 28132 19796 28138 19848
rect 28184 19836 28212 19876
rect 29086 19864 29092 19916
rect 29144 19904 29150 19916
rect 29181 19907 29239 19913
rect 29181 19904 29193 19907
rect 29144 19876 29193 19904
rect 29144 19864 29150 19876
rect 29181 19873 29193 19876
rect 29227 19873 29239 19907
rect 29181 19867 29239 19873
rect 29270 19864 29276 19916
rect 29328 19904 29334 19916
rect 30009 19907 30067 19913
rect 30009 19904 30021 19907
rect 29328 19876 30021 19904
rect 29328 19864 29334 19876
rect 30009 19873 30021 19876
rect 30055 19873 30067 19907
rect 30009 19867 30067 19873
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 28184 19808 29745 19836
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 30374 19796 30380 19848
rect 30432 19836 30438 19848
rect 31404 19836 31432 20012
rect 34330 20000 34336 20052
rect 34388 20040 34394 20052
rect 34701 20043 34759 20049
rect 34701 20040 34713 20043
rect 34388 20012 34713 20040
rect 34388 20000 34394 20012
rect 34701 20009 34713 20012
rect 34747 20009 34759 20043
rect 34701 20003 34759 20009
rect 31478 19864 31484 19916
rect 31536 19904 31542 19916
rect 31573 19907 31631 19913
rect 31573 19904 31585 19907
rect 31536 19876 31585 19904
rect 31536 19864 31542 19876
rect 31573 19873 31585 19876
rect 31619 19873 31631 19907
rect 31573 19867 31631 19873
rect 31662 19864 31668 19916
rect 31720 19904 31726 19916
rect 33505 19907 33563 19913
rect 33505 19904 33517 19907
rect 31720 19876 33517 19904
rect 31720 19864 31726 19876
rect 33505 19873 33517 19876
rect 33551 19873 33563 19907
rect 33505 19867 33563 19873
rect 33594 19864 33600 19916
rect 33652 19904 33658 19916
rect 33781 19907 33839 19913
rect 33781 19904 33793 19907
rect 33652 19876 33793 19904
rect 33652 19864 33658 19876
rect 33781 19873 33793 19876
rect 33827 19873 33839 19907
rect 33781 19867 33839 19873
rect 32217 19839 32275 19845
rect 32217 19836 32229 19839
rect 30432 19808 31156 19836
rect 31404 19808 32229 19836
rect 30432 19796 30438 19808
rect 26142 19768 26148 19780
rect 25332 19740 26148 19768
rect 26142 19728 26148 19740
rect 26200 19728 26206 19780
rect 26878 19728 26884 19780
rect 26936 19728 26942 19780
rect 31128 19768 31156 19808
rect 32217 19805 32229 19808
rect 32263 19836 32275 19839
rect 33137 19839 33195 19845
rect 33137 19836 33149 19839
rect 32263 19808 33149 19836
rect 32263 19805 32275 19808
rect 32217 19799 32275 19805
rect 33137 19805 33149 19808
rect 33183 19805 33195 19839
rect 33137 19799 33195 19805
rect 31386 19768 31392 19780
rect 27540 19740 31064 19768
rect 31128 19740 31392 19768
rect 24673 19703 24731 19709
rect 24673 19669 24685 19703
rect 24719 19669 24731 19703
rect 24673 19663 24731 19669
rect 25133 19703 25191 19709
rect 25133 19669 25145 19703
rect 25179 19700 25191 19703
rect 27540 19700 27568 19740
rect 25179 19672 27568 19700
rect 25179 19669 25191 19672
rect 25133 19663 25191 19669
rect 28718 19660 28724 19712
rect 28776 19660 28782 19712
rect 29089 19703 29147 19709
rect 29089 19669 29101 19703
rect 29135 19700 29147 19703
rect 29362 19700 29368 19712
rect 29135 19672 29368 19700
rect 29135 19669 29147 19672
rect 29089 19663 29147 19669
rect 29362 19660 29368 19672
rect 29420 19660 29426 19712
rect 31036 19709 31064 19740
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 31481 19771 31539 19777
rect 31481 19737 31493 19771
rect 31527 19768 31539 19771
rect 41966 19768 41972 19780
rect 31527 19740 41972 19768
rect 31527 19737 31539 19740
rect 31481 19731 31539 19737
rect 41966 19728 41972 19740
rect 42024 19728 42030 19780
rect 31021 19703 31079 19709
rect 31021 19669 31033 19703
rect 31067 19669 31079 19703
rect 31021 19663 31079 19669
rect 31570 19660 31576 19712
rect 31628 19700 31634 19712
rect 32861 19703 32919 19709
rect 32861 19700 32873 19703
rect 31628 19672 32873 19700
rect 31628 19660 31634 19672
rect 32861 19669 32873 19672
rect 32907 19669 32919 19703
rect 32861 19663 32919 19669
rect 34882 19660 34888 19712
rect 34940 19660 34946 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 3605 19499 3663 19505
rect 3605 19496 3617 19499
rect 1820 19468 3617 19496
rect 1820 19456 1826 19468
rect 3605 19465 3617 19468
rect 3651 19465 3663 19499
rect 3605 19459 3663 19465
rect 3786 19456 3792 19508
rect 3844 19496 3850 19508
rect 4522 19496 4528 19508
rect 3844 19468 4528 19496
rect 3844 19456 3850 19468
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 4890 19456 4896 19508
rect 4948 19456 4954 19508
rect 5997 19499 6055 19505
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 6086 19496 6092 19508
rect 6043 19468 6092 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 6270 19456 6276 19508
rect 6328 19496 6334 19508
rect 6638 19496 6644 19508
rect 6328 19468 6644 19496
rect 6328 19456 6334 19468
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 9033 19499 9091 19505
rect 9033 19496 9045 19499
rect 8996 19468 9045 19496
rect 8996 19456 9002 19468
rect 9033 19465 9045 19468
rect 9079 19465 9091 19499
rect 9033 19459 9091 19465
rect 9766 19456 9772 19508
rect 9824 19456 9830 19508
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 10008 19468 10241 19496
rect 10008 19456 10014 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 11164 19468 13308 19496
rect 3694 19428 3700 19440
rect 1780 19400 3700 19428
rect 1780 19369 1808 19400
rect 3694 19388 3700 19400
rect 3752 19388 3758 19440
rect 4908 19428 4936 19456
rect 4264 19400 4936 19428
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19329 1823 19363
rect 1765 19323 1823 19329
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 4264 19369 4292 19400
rect 5810 19388 5816 19440
rect 5868 19428 5874 19440
rect 7466 19428 7472 19440
rect 5868 19400 7472 19428
rect 5868 19388 5874 19400
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 7616 19400 8050 19428
rect 7616 19388 7622 19400
rect 9122 19388 9128 19440
rect 9180 19428 9186 19440
rect 11054 19428 11060 19440
rect 9180 19400 11060 19428
rect 9180 19388 9186 19400
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 3789 19363 3847 19369
rect 3789 19360 3801 19363
rect 3660 19332 3801 19360
rect 3660 19320 3666 19332
rect 3789 19329 3801 19332
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 6270 19360 6276 19372
rect 5684 19332 6276 19360
rect 5684 19320 5690 19332
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 7282 19360 7288 19372
rect 6880 19332 7288 19360
rect 6880 19320 6886 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 10134 19360 10140 19372
rect 9723 19332 10140 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 11164 19369 11192 19468
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 11480 19400 12466 19428
rect 11480 19388 11486 19400
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 13280 19360 13308 19468
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 14056 19468 17877 19496
rect 14056 19456 14062 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 18322 19456 18328 19508
rect 18380 19456 18386 19508
rect 18506 19456 18512 19508
rect 18564 19496 18570 19508
rect 19061 19499 19119 19505
rect 19061 19496 19073 19499
rect 18564 19468 19073 19496
rect 18564 19456 18570 19468
rect 19061 19465 19073 19468
rect 19107 19465 19119 19499
rect 19061 19459 19119 19465
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 20622 19496 20628 19508
rect 19300 19468 20628 19496
rect 19300 19456 19306 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21453 19499 21511 19505
rect 21453 19496 21465 19499
rect 20864 19468 21465 19496
rect 20864 19456 20870 19468
rect 21453 19465 21465 19468
rect 21499 19496 21511 19499
rect 21499 19468 22094 19496
rect 21499 19465 21511 19468
rect 21453 19459 21511 19465
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 14645 19431 14703 19437
rect 14645 19428 14657 19431
rect 13780 19400 14657 19428
rect 13780 19388 13786 19400
rect 14645 19397 14657 19400
rect 14691 19397 14703 19431
rect 14645 19391 14703 19397
rect 15010 19388 15016 19440
rect 15068 19428 15074 19440
rect 15068 19400 17632 19428
rect 15068 19388 15074 19400
rect 13814 19360 13820 19372
rect 13280 19332 13820 19360
rect 13814 19320 13820 19332
rect 13872 19320 13878 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19329 13967 19363
rect 13909 19323 13967 19329
rect 4522 19252 4528 19304
rect 4580 19252 4586 19304
rect 5074 19252 5080 19304
rect 5132 19292 5138 19304
rect 5644 19292 5672 19320
rect 5132 19264 5672 19292
rect 5132 19252 5138 19264
rect 5810 19252 5816 19304
rect 5868 19292 5874 19304
rect 7561 19295 7619 19301
rect 7561 19292 7573 19295
rect 5868 19264 7573 19292
rect 5868 19252 5874 19264
rect 7561 19261 7573 19264
rect 7607 19261 7619 19295
rect 7561 19255 7619 19261
rect 10410 19252 10416 19304
rect 10468 19252 10474 19304
rect 10502 19252 10508 19304
rect 10560 19292 10566 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 10560 19264 11989 19292
rect 10560 19252 10566 19264
rect 11977 19261 11989 19264
rect 12023 19292 12035 19295
rect 12066 19292 12072 19304
rect 12023 19264 12072 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 12676 19264 13461 19292
rect 12676 19252 12682 19264
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13924 19292 13952 19323
rect 14274 19320 14280 19372
rect 14332 19360 14338 19372
rect 14734 19360 14740 19372
rect 14332 19332 14740 19360
rect 14332 19320 14338 19332
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16574 19360 16580 19372
rect 15804 19332 16580 19360
rect 15804 19320 15810 19332
rect 16574 19320 16580 19332
rect 16632 19320 16638 19372
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17310 19360 17316 19372
rect 16991 19332 17316 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 13998 19292 14004 19304
rect 13924 19264 14004 19292
rect 3326 19184 3332 19236
rect 3384 19184 3390 19236
rect 6825 19227 6883 19233
rect 6825 19224 6837 19227
rect 5552 19196 6837 19224
rect 3786 19116 3792 19168
rect 3844 19156 3850 19168
rect 5552 19156 5580 19196
rect 6825 19193 6837 19196
rect 6871 19193 6883 19227
rect 13924 19224 13952 19264
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 14148 19264 15853 19292
rect 14148 19252 14154 19264
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 17218 19292 17224 19304
rect 15841 19255 15899 19261
rect 16132 19264 17224 19292
rect 6825 19187 6883 19193
rect 9416 19196 11836 19224
rect 3844 19128 5580 19156
rect 3844 19116 3850 19128
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 6914 19156 6920 19168
rect 6328 19128 6920 19156
rect 6328 19116 6334 19128
rect 6914 19116 6920 19128
rect 6972 19156 6978 19168
rect 7558 19156 7564 19168
rect 6972 19128 7564 19156
rect 6972 19116 6978 19128
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 9416 19165 9444 19196
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 9180 19128 9413 19156
rect 9180 19116 9186 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10836 19128 10977 19156
rect 10836 19116 10842 19128
rect 10965 19125 10977 19128
rect 11011 19125 11023 19159
rect 10965 19119 11023 19125
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11422 19156 11428 19168
rect 11204 19128 11428 19156
rect 11204 19116 11210 19128
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 11808 19156 11836 19196
rect 13004 19196 13952 19224
rect 13004 19156 13032 19196
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14240 19196 15301 19224
rect 14240 19184 14246 19196
rect 15289 19193 15301 19196
rect 15335 19193 15347 19227
rect 15289 19187 15347 19193
rect 11808 19128 13032 19156
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13538 19156 13544 19168
rect 13136 19128 13544 19156
rect 13136 19116 13142 19128
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 15010 19156 15016 19168
rect 13780 19128 15016 19156
rect 13780 19116 13786 19128
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 16132 19156 16160 19264
rect 17218 19252 17224 19264
rect 17276 19292 17282 19304
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 17276 19264 17509 19292
rect 17276 19252 17282 19264
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17604 19292 17632 19400
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 20254 19428 20260 19440
rect 19392 19400 20260 19428
rect 19392 19388 19398 19400
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 20530 19388 20536 19440
rect 20588 19388 20594 19440
rect 22066 19428 22094 19468
rect 22462 19456 22468 19508
rect 22520 19456 22526 19508
rect 22830 19456 22836 19508
rect 22888 19456 22894 19508
rect 22925 19499 22983 19505
rect 22925 19465 22937 19499
rect 22971 19496 22983 19499
rect 23842 19496 23848 19508
rect 22971 19468 23848 19496
rect 22971 19465 22983 19468
rect 22925 19459 22983 19465
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 24121 19499 24179 19505
rect 24121 19465 24133 19499
rect 24167 19496 24179 19499
rect 26234 19496 26240 19508
rect 24167 19468 26240 19496
rect 24167 19465 24179 19468
rect 24121 19459 24179 19465
rect 26234 19456 26240 19468
rect 26292 19456 26298 19508
rect 26326 19456 26332 19508
rect 26384 19496 26390 19508
rect 30101 19499 30159 19505
rect 26384 19468 29960 19496
rect 26384 19456 26390 19468
rect 23750 19428 23756 19440
rect 22066 19400 23756 19428
rect 23750 19388 23756 19400
rect 23808 19428 23814 19440
rect 23808 19400 24256 19428
rect 23808 19388 23814 19400
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18598 19320 18604 19372
rect 18656 19320 18662 19372
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 17604 19264 18429 19292
rect 17497 19255 17555 19261
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 16206 19184 16212 19236
rect 16264 19224 16270 19236
rect 18616 19224 18644 19320
rect 19702 19292 19708 19304
rect 19306 19264 19708 19292
rect 19306 19224 19334 19264
rect 19702 19252 19708 19264
rect 19760 19252 19766 19304
rect 19978 19252 19984 19304
rect 20036 19252 20042 19304
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20622 19292 20628 19304
rect 20128 19264 20628 19292
rect 20128 19252 20134 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21910 19292 21916 19304
rect 20772 19264 21916 19292
rect 20772 19252 20778 19264
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 24228 19301 24256 19400
rect 25774 19388 25780 19440
rect 25832 19388 25838 19440
rect 28902 19428 28908 19440
rect 26436 19400 28908 19428
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 25038 19360 25044 19372
rect 24995 19332 25044 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19292 23167 19295
rect 24213 19295 24271 19301
rect 23155 19264 23888 19292
rect 23155 19261 23167 19264
rect 23109 19255 23167 19261
rect 23661 19227 23719 19233
rect 23661 19224 23673 19227
rect 16264 19196 19334 19224
rect 21008 19196 23673 19224
rect 16264 19184 16270 19196
rect 15252 19128 16160 19156
rect 15252 19116 15258 19128
rect 16482 19116 16488 19168
rect 16540 19116 16546 19168
rect 16850 19116 16856 19168
rect 16908 19156 16914 19168
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 16908 19128 17049 19156
rect 16908 19116 16914 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 21008 19156 21036 19196
rect 23661 19193 23673 19196
rect 23707 19193 23719 19227
rect 23661 19187 23719 19193
rect 18564 19128 21036 19156
rect 18564 19116 18570 19128
rect 22186 19116 22192 19168
rect 22244 19116 22250 19168
rect 23860 19156 23888 19264
rect 24213 19261 24225 19295
rect 24259 19261 24271 19295
rect 24213 19255 24271 19261
rect 23934 19184 23940 19236
rect 23992 19224 23998 19236
rect 26436 19233 26464 19400
rect 28902 19388 28908 19400
rect 28960 19388 28966 19440
rect 29362 19388 29368 19440
rect 29420 19388 29426 19440
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 26605 19363 26663 19369
rect 26605 19360 26617 19363
rect 26568 19332 26617 19360
rect 26568 19320 26574 19332
rect 26605 19329 26617 19332
rect 26651 19329 26663 19363
rect 26605 19323 26663 19329
rect 27246 19320 27252 19372
rect 27304 19320 27310 19372
rect 27798 19320 27804 19372
rect 27856 19360 27862 19372
rect 27893 19363 27951 19369
rect 27893 19360 27905 19363
rect 27856 19332 27905 19360
rect 27856 19320 27862 19332
rect 27893 19329 27905 19332
rect 27939 19329 27951 19363
rect 27893 19323 27951 19329
rect 28350 19320 28356 19372
rect 28408 19320 28414 19372
rect 29932 19360 29960 19468
rect 30101 19465 30113 19499
rect 30147 19496 30159 19499
rect 31202 19496 31208 19508
rect 30147 19468 31208 19496
rect 30147 19465 30159 19468
rect 30101 19459 30159 19465
rect 31202 19456 31208 19468
rect 31260 19456 31266 19508
rect 31294 19456 31300 19508
rect 31352 19496 31358 19508
rect 37550 19496 37556 19508
rect 31352 19468 37556 19496
rect 31352 19456 31358 19468
rect 37550 19456 37556 19468
rect 37608 19456 37614 19508
rect 31386 19388 31392 19440
rect 31444 19428 31450 19440
rect 31665 19431 31723 19437
rect 31665 19428 31677 19431
rect 31444 19400 31677 19428
rect 31444 19388 31450 19400
rect 31665 19397 31677 19400
rect 31711 19428 31723 19431
rect 31846 19428 31852 19440
rect 31711 19400 31852 19428
rect 31711 19397 31723 19400
rect 31665 19391 31723 19397
rect 31846 19388 31852 19400
rect 31904 19388 31910 19440
rect 32398 19388 32404 19440
rect 32456 19388 32462 19440
rect 33134 19388 33140 19440
rect 33192 19428 33198 19440
rect 33597 19431 33655 19437
rect 33597 19428 33609 19431
rect 33192 19400 33609 19428
rect 33192 19388 33198 19400
rect 33597 19397 33609 19400
rect 33643 19397 33655 19431
rect 33597 19391 33655 19397
rect 30561 19363 30619 19369
rect 30561 19360 30573 19363
rect 29932 19332 30573 19360
rect 30561 19329 30573 19332
rect 30607 19329 30619 19363
rect 30561 19323 30619 19329
rect 30650 19320 30656 19372
rect 30708 19360 30714 19372
rect 31205 19363 31263 19369
rect 31205 19360 31217 19363
rect 30708 19332 31217 19360
rect 30708 19320 30714 19332
rect 31205 19329 31217 19332
rect 31251 19329 31263 19363
rect 31754 19360 31760 19372
rect 31205 19323 31263 19329
rect 31680 19332 31760 19360
rect 28629 19295 28687 19301
rect 28629 19261 28641 19295
rect 28675 19292 28687 19295
rect 29178 19292 29184 19304
rect 28675 19264 29184 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 29178 19252 29184 19264
rect 29236 19252 29242 19304
rect 29362 19252 29368 19304
rect 29420 19292 29426 19304
rect 29822 19292 29828 19304
rect 29420 19264 29828 19292
rect 29420 19252 29426 19264
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 31573 19295 31631 19301
rect 31573 19261 31585 19295
rect 31619 19292 31631 19295
rect 31680 19292 31708 19332
rect 31754 19320 31760 19332
rect 31812 19320 31818 19372
rect 31619 19264 31708 19292
rect 31941 19295 31999 19301
rect 31619 19261 31631 19264
rect 31573 19255 31631 19261
rect 31941 19261 31953 19295
rect 31987 19292 31999 19295
rect 32306 19292 32312 19304
rect 31987 19264 32312 19292
rect 31987 19261 31999 19264
rect 31941 19255 31999 19261
rect 32306 19252 32312 19264
rect 32364 19252 32370 19304
rect 32398 19252 32404 19304
rect 32456 19292 32462 19304
rect 39758 19292 39764 19304
rect 32456 19264 39764 19292
rect 32456 19252 32462 19264
rect 39758 19252 39764 19264
rect 39816 19252 39822 19304
rect 26421 19227 26479 19233
rect 23992 19196 26372 19224
rect 23992 19184 23998 19196
rect 26142 19156 26148 19168
rect 23860 19128 26148 19156
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 26234 19116 26240 19168
rect 26292 19116 26298 19168
rect 26344 19156 26372 19196
rect 26421 19193 26433 19227
rect 26467 19193 26479 19227
rect 45830 19224 45836 19236
rect 26421 19187 26479 19193
rect 29656 19196 45836 19224
rect 29656 19156 29684 19196
rect 45830 19184 45836 19196
rect 45888 19184 45894 19236
rect 26344 19128 29684 19156
rect 32490 19116 32496 19168
rect 32548 19116 32554 19168
rect 33229 19159 33287 19165
rect 33229 19125 33241 19159
rect 33275 19156 33287 19159
rect 33318 19156 33324 19168
rect 33275 19128 33324 19156
rect 33275 19125 33287 19128
rect 33229 19119 33287 19125
rect 33318 19116 33324 19128
rect 33376 19116 33382 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 3418 18912 3424 18964
rect 3476 18952 3482 18964
rect 3881 18955 3939 18961
rect 3881 18952 3893 18955
rect 3476 18924 3893 18952
rect 3476 18912 3482 18924
rect 3881 18921 3893 18924
rect 3927 18952 3939 18955
rect 9122 18952 9128 18964
rect 3927 18924 9128 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 10410 18912 10416 18964
rect 10468 18952 10474 18964
rect 12434 18952 12440 18964
rect 10468 18924 12440 18952
rect 10468 18912 10474 18924
rect 12434 18912 12440 18924
rect 12492 18952 12498 18964
rect 13722 18952 13728 18964
rect 12492 18924 13728 18952
rect 12492 18912 12498 18924
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14277 18955 14335 18961
rect 14277 18921 14289 18955
rect 14323 18952 14335 18955
rect 14458 18952 14464 18964
rect 14323 18924 14464 18952
rect 14323 18921 14335 18924
rect 14277 18915 14335 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 15120 18924 18153 18952
rect 3602 18844 3608 18896
rect 3660 18844 3666 18896
rect 4065 18887 4123 18893
rect 4065 18853 4077 18887
rect 4111 18884 4123 18887
rect 5074 18884 5080 18896
rect 4111 18856 5080 18884
rect 4111 18853 4123 18856
rect 4065 18847 4123 18853
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 10594 18844 10600 18896
rect 10652 18844 10658 18896
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 11020 18856 11376 18884
rect 11020 18844 11026 18856
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1452 18788 2053 18816
rect 1452 18776 1458 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18816 3479 18819
rect 4154 18816 4160 18828
rect 3467 18788 4160 18816
rect 3467 18785 3479 18788
rect 3421 18779 3479 18785
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5350 18816 5356 18828
rect 5031 18788 5356 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18816 5595 18819
rect 6822 18816 6828 18828
rect 5583 18788 6828 18816
rect 5583 18785 5595 18788
rect 5537 18779 5595 18785
rect 6822 18776 6828 18788
rect 6880 18776 6886 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7834 18816 7840 18828
rect 7432 18788 7840 18816
rect 7432 18776 7438 18788
rect 7834 18776 7840 18788
rect 7892 18816 7898 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 7892 18788 8401 18816
rect 7892 18776 7898 18788
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 8628 18788 9781 18816
rect 8628 18776 8634 18788
rect 9769 18785 9781 18788
rect 9815 18785 9827 18819
rect 9769 18779 9827 18785
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10318 18816 10324 18828
rect 10192 18788 10324 18816
rect 10192 18776 10198 18788
rect 10318 18776 10324 18788
rect 10376 18776 10382 18828
rect 10686 18776 10692 18828
rect 10744 18816 10750 18828
rect 10870 18816 10876 18828
rect 10744 18788 10876 18816
rect 10744 18776 10750 18788
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18785 11299 18819
rect 11241 18779 11299 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 1854 18748 1860 18760
rect 1811 18720 1860 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 1854 18708 1860 18720
rect 1912 18708 1918 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4755 18720 5580 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 5258 18680 5264 18692
rect 4356 18652 5264 18680
rect 4356 18621 4384 18652
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 4341 18615 4399 18621
rect 4341 18581 4353 18615
rect 4387 18581 4399 18615
rect 4341 18575 4399 18581
rect 4798 18572 4804 18624
rect 4856 18572 4862 18624
rect 5552 18612 5580 18720
rect 6914 18708 6920 18760
rect 6972 18708 6978 18760
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18748 7803 18751
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 7791 18720 8217 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 8205 18717 8217 18720
rect 8251 18748 8263 18751
rect 8294 18748 8300 18760
rect 8251 18720 8300 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18748 9643 18751
rect 10410 18748 10416 18760
rect 9631 18720 10416 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10965 18751 11023 18757
rect 10965 18744 10977 18751
rect 10888 18717 10977 18744
rect 11011 18717 11023 18751
rect 10888 18716 11023 18717
rect 5813 18683 5871 18689
rect 5813 18649 5825 18683
rect 5859 18680 5871 18683
rect 5902 18680 5908 18692
rect 5859 18652 5908 18680
rect 5859 18649 5871 18652
rect 5813 18643 5871 18649
rect 5902 18640 5908 18652
rect 5960 18640 5966 18692
rect 8386 18680 8392 18692
rect 7208 18652 8392 18680
rect 7208 18612 7236 18652
rect 8386 18640 8392 18652
rect 8444 18680 8450 18692
rect 9398 18680 9404 18692
rect 8444 18652 9404 18680
rect 8444 18640 8450 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 10505 18683 10563 18689
rect 10505 18680 10517 18683
rect 9824 18652 10517 18680
rect 9824 18640 9830 18652
rect 10505 18649 10517 18652
rect 10551 18680 10563 18683
rect 10888 18680 10916 18716
rect 10965 18711 11023 18716
rect 10551 18652 10916 18680
rect 10551 18649 10563 18652
rect 10505 18643 10563 18649
rect 11256 18624 11284 18779
rect 11348 18748 11376 18856
rect 11606 18844 11612 18896
rect 11664 18884 11670 18896
rect 11793 18887 11851 18893
rect 11793 18884 11805 18887
rect 11664 18856 11805 18884
rect 11664 18844 11670 18856
rect 11793 18853 11805 18856
rect 11839 18853 11851 18887
rect 11793 18847 11851 18853
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 14553 18887 14611 18893
rect 14553 18884 14565 18887
rect 12584 18856 14565 18884
rect 12584 18844 12590 18856
rect 14553 18853 14565 18856
rect 14599 18853 14611 18887
rect 14553 18847 14611 18853
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12216 18788 12357 18816
rect 12216 18776 12222 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 15010 18816 15016 18828
rect 12345 18779 12403 18785
rect 13096 18788 15016 18816
rect 11348 18720 11928 18748
rect 11701 18683 11759 18689
rect 11701 18649 11713 18683
rect 11747 18680 11759 18683
rect 11790 18680 11796 18692
rect 11747 18652 11796 18680
rect 11747 18649 11759 18652
rect 11701 18643 11759 18649
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 11900 18680 11928 18720
rect 11974 18708 11980 18760
rect 12032 18748 12038 18760
rect 12618 18748 12624 18760
rect 12032 18720 12624 18748
rect 12032 18708 12038 18720
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 13096 18757 13124 18788
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 13069 18751 13127 18757
rect 13069 18717 13081 18751
rect 13115 18717 13127 18751
rect 13069 18711 13127 18717
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 15120 18748 15148 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 19242 18952 19248 18964
rect 18141 18915 18199 18921
rect 18524 18924 19248 18952
rect 16758 18844 16764 18896
rect 16816 18884 16822 18896
rect 17681 18887 17739 18893
rect 17681 18884 17693 18887
rect 16816 18856 17693 18884
rect 16816 18844 16822 18856
rect 17681 18853 17693 18856
rect 17727 18853 17739 18887
rect 17681 18847 17739 18853
rect 17770 18844 17776 18896
rect 17828 18884 17834 18896
rect 18524 18884 18552 18924
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19334 18912 19340 18964
rect 19392 18912 19398 18964
rect 20070 18952 20076 18964
rect 19444 18924 20076 18952
rect 17828 18856 18552 18884
rect 17828 18844 17834 18856
rect 18598 18844 18604 18896
rect 18656 18884 18662 18896
rect 19444 18884 19472 18924
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 22186 18952 22192 18964
rect 20272 18924 22192 18952
rect 20272 18884 20300 18924
rect 22186 18912 22192 18924
rect 22244 18952 22250 18964
rect 23382 18952 23388 18964
rect 22244 18924 23388 18952
rect 22244 18912 22250 18924
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 25672 18955 25730 18961
rect 25672 18921 25684 18955
rect 25718 18952 25730 18955
rect 28718 18952 28724 18964
rect 25718 18924 28724 18952
rect 25718 18921 25730 18924
rect 25672 18915 25730 18921
rect 28718 18912 28724 18924
rect 28776 18912 28782 18964
rect 28810 18912 28816 18964
rect 28868 18912 28874 18964
rect 28994 18912 29000 18964
rect 29052 18952 29058 18964
rect 32953 18955 33011 18961
rect 32953 18952 32965 18955
rect 29052 18924 32965 18952
rect 29052 18912 29058 18924
rect 28442 18884 28448 18896
rect 18656 18856 19472 18884
rect 20088 18856 20300 18884
rect 27172 18856 28448 18884
rect 18656 18844 18662 18856
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 16206 18816 16212 18828
rect 15243 18788 16212 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 16206 18776 16212 18788
rect 16264 18776 16270 18828
rect 16942 18816 16948 18828
rect 16500 18788 16948 18816
rect 14783 18720 15148 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 16500 18692 16528 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 18690 18816 18696 18828
rect 17184 18788 18696 18816
rect 17184 18776 17190 18788
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 20088 18816 20116 18856
rect 19628 18788 20116 18816
rect 16776 18720 17632 18748
rect 14274 18680 14280 18692
rect 11900 18652 14280 18680
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 16482 18640 16488 18692
rect 16540 18640 16546 18692
rect 5552 18584 7236 18612
rect 7282 18572 7288 18624
rect 7340 18572 7346 18624
rect 7834 18572 7840 18624
rect 7892 18572 7898 18624
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 9030 18612 9036 18624
rect 8343 18584 9036 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9214 18572 9220 18624
rect 9272 18572 9278 18624
rect 9490 18572 9496 18624
rect 9548 18612 9554 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9548 18584 9689 18612
rect 9548 18572 9554 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9677 18575 9735 18581
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 11054 18572 11060 18624
rect 11112 18572 11118 18624
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11974 18612 11980 18624
rect 11296 18584 11980 18612
rect 11296 18572 11302 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12161 18615 12219 18621
rect 12161 18612 12173 18615
rect 12124 18584 12173 18612
rect 12124 18572 12130 18584
rect 12161 18581 12173 18584
rect 12207 18581 12219 18615
rect 12161 18575 12219 18581
rect 12250 18572 12256 18624
rect 12308 18572 12314 18624
rect 13725 18615 13783 18621
rect 13725 18581 13737 18615
rect 13771 18612 13783 18615
rect 16776 18612 16804 18720
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 17497 18683 17555 18689
rect 17497 18680 17509 18683
rect 17276 18652 17509 18680
rect 17276 18640 17282 18652
rect 17497 18649 17509 18652
rect 17543 18649 17555 18683
rect 17604 18680 17632 18720
rect 18506 18708 18512 18760
rect 18564 18708 18570 18760
rect 19628 18757 19656 18788
rect 20162 18776 20168 18828
rect 20220 18816 20226 18828
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20220 18788 21189 18816
rect 20220 18776 20226 18788
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 21450 18776 21456 18828
rect 21508 18776 21514 18828
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 23934 18816 23940 18828
rect 21876 18788 23940 18816
rect 21876 18776 21882 18788
rect 23934 18776 23940 18788
rect 23992 18776 23998 18828
rect 24026 18776 24032 18828
rect 24084 18816 24090 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24084 18788 24593 18816
rect 24084 18776 24090 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25774 18816 25780 18828
rect 25455 18788 25780 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 26142 18776 26148 18828
rect 26200 18816 26206 18828
rect 27172 18825 27200 18856
rect 28442 18844 28448 18856
rect 28500 18844 28506 18896
rect 28626 18844 28632 18896
rect 28684 18844 28690 18896
rect 32398 18884 32404 18896
rect 30300 18856 32404 18884
rect 27157 18819 27215 18825
rect 27157 18816 27169 18819
rect 26200 18788 27169 18816
rect 26200 18776 26206 18788
rect 27157 18785 27169 18788
rect 27203 18785 27215 18819
rect 27157 18779 27215 18785
rect 27246 18776 27252 18828
rect 27304 18816 27310 18828
rect 28261 18819 28319 18825
rect 28261 18816 28273 18819
rect 27304 18788 28273 18816
rect 27304 18776 27310 18788
rect 28261 18785 28273 18788
rect 28307 18816 28319 18819
rect 29822 18816 29828 18828
rect 28307 18788 29828 18816
rect 28307 18785 28319 18788
rect 28261 18779 28319 18785
rect 29822 18776 29828 18788
rect 29880 18776 29886 18828
rect 30006 18776 30012 18828
rect 30064 18816 30070 18828
rect 30300 18825 30328 18856
rect 32398 18844 32404 18856
rect 32456 18844 32462 18896
rect 32493 18887 32551 18893
rect 32493 18853 32505 18887
rect 32539 18884 32551 18887
rect 32582 18884 32588 18896
rect 32539 18856 32588 18884
rect 32539 18853 32551 18856
rect 32493 18847 32551 18853
rect 32582 18844 32588 18856
rect 32640 18844 32646 18896
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 30064 18788 30297 18816
rect 30064 18776 30070 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 32122 18816 32128 18828
rect 30285 18779 30343 18785
rect 30852 18788 32128 18816
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 19760 18720 20361 18748
rect 19760 18708 19766 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22520 18720 22586 18748
rect 22520 18708 22526 18720
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 23385 18751 23443 18757
rect 23385 18748 23397 18751
rect 23348 18720 23397 18748
rect 23348 18708 23354 18720
rect 23385 18717 23397 18720
rect 23431 18717 23443 18751
rect 23385 18711 23443 18717
rect 26786 18708 26792 18760
rect 26844 18708 26850 18760
rect 28626 18708 28632 18760
rect 28684 18748 28690 18760
rect 28997 18751 29055 18757
rect 28997 18748 29009 18751
rect 28684 18720 29009 18748
rect 28684 18708 28690 18720
rect 28997 18717 29009 18720
rect 29043 18717 29055 18751
rect 28997 18711 29055 18717
rect 30190 18708 30196 18760
rect 30248 18748 30254 18760
rect 30852 18748 30880 18788
rect 32122 18776 32128 18788
rect 32180 18776 32186 18828
rect 30248 18720 30880 18748
rect 30929 18751 30987 18757
rect 30248 18708 30254 18720
rect 30929 18717 30941 18751
rect 30975 18748 30987 18751
rect 31202 18748 31208 18760
rect 30975 18720 31208 18748
rect 30975 18717 30987 18720
rect 30929 18711 30987 18717
rect 31202 18708 31208 18720
rect 31260 18708 31266 18760
rect 32677 18751 32735 18757
rect 32677 18717 32689 18751
rect 32723 18748 32735 18751
rect 32784 18748 32812 18924
rect 32953 18921 32965 18924
rect 32999 18921 33011 18955
rect 32953 18915 33011 18921
rect 32723 18720 32812 18748
rect 32723 18717 32735 18720
rect 32677 18711 32735 18717
rect 19978 18680 19984 18692
rect 17604 18652 19984 18680
rect 17497 18643 17555 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 20088 18652 20944 18680
rect 22678 18652 23152 18680
rect 13771 18584 16804 18612
rect 13771 18581 13783 18584
rect 13725 18575 13783 18581
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17402 18612 17408 18624
rect 17000 18584 17408 18612
rect 17000 18572 17006 18584
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18506 18612 18512 18624
rect 18288 18584 18512 18612
rect 18288 18572 18294 18584
rect 18506 18572 18512 18584
rect 18564 18572 18570 18624
rect 18598 18572 18604 18624
rect 18656 18572 18662 18624
rect 18690 18572 18696 18624
rect 18748 18612 18754 18624
rect 20088 18612 20116 18652
rect 18748 18584 20116 18612
rect 18748 18572 18754 18584
rect 20806 18572 20812 18624
rect 20864 18572 20870 18624
rect 20916 18612 20944 18652
rect 22925 18615 22983 18621
rect 22925 18612 22937 18615
rect 20916 18584 22937 18612
rect 22925 18581 22937 18584
rect 22971 18581 22983 18615
rect 23124 18612 23152 18652
rect 23198 18640 23204 18692
rect 23256 18680 23262 18692
rect 25958 18680 25964 18692
rect 23256 18652 25964 18680
rect 23256 18640 23262 18652
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 28077 18683 28135 18689
rect 28077 18649 28089 18683
rect 28123 18680 28135 18683
rect 29914 18680 29920 18692
rect 28123 18652 29920 18680
rect 28123 18649 28135 18652
rect 28077 18643 28135 18649
rect 29914 18640 29920 18652
rect 29972 18640 29978 18692
rect 30098 18640 30104 18692
rect 30156 18680 30162 18692
rect 31941 18683 31999 18689
rect 31941 18680 31953 18683
rect 30156 18652 31953 18680
rect 30156 18640 30162 18652
rect 31941 18649 31953 18652
rect 31987 18680 31999 18683
rect 42518 18680 42524 18692
rect 31987 18652 42524 18680
rect 31987 18649 31999 18652
rect 31941 18643 31999 18649
rect 42518 18640 42524 18652
rect 42576 18640 42582 18692
rect 23842 18612 23848 18624
rect 23124 18584 23848 18612
rect 22925 18575 22983 18581
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 24029 18615 24087 18621
rect 24029 18581 24041 18615
rect 24075 18612 24087 18615
rect 24854 18612 24860 18624
rect 24075 18584 24860 18612
rect 24075 18581 24087 18584
rect 24029 18575 24087 18581
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 25038 18572 25044 18624
rect 25096 18572 25102 18624
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 27617 18615 27675 18621
rect 27617 18612 27629 18615
rect 25188 18584 27629 18612
rect 25188 18572 25194 18584
rect 27617 18581 27629 18584
rect 27663 18581 27675 18615
rect 27617 18575 27675 18581
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 27985 18615 28043 18621
rect 27985 18612 27997 18615
rect 27764 18584 27997 18612
rect 27764 18572 27770 18584
rect 27985 18581 27997 18584
rect 28031 18581 28043 18615
rect 27985 18575 28043 18581
rect 29365 18615 29423 18621
rect 29365 18581 29377 18615
rect 29411 18612 29423 18615
rect 29454 18612 29460 18624
rect 29411 18584 29460 18612
rect 29411 18581 29423 18584
rect 29365 18575 29423 18581
rect 29454 18572 29460 18584
rect 29512 18572 29518 18624
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30282 18572 30288 18624
rect 30340 18612 30346 18624
rect 31573 18615 31631 18621
rect 31573 18612 31585 18615
rect 30340 18584 31585 18612
rect 30340 18572 30346 18584
rect 31573 18581 31585 18584
rect 31619 18581 31631 18615
rect 31573 18575 31631 18581
rect 32122 18572 32128 18624
rect 32180 18612 32186 18624
rect 43714 18612 43720 18624
rect 32180 18584 43720 18612
rect 32180 18572 32186 18584
rect 43714 18572 43720 18584
rect 43772 18572 43778 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 2280 18380 3924 18408
rect 2280 18368 2286 18380
rect 3786 18340 3792 18352
rect 1780 18312 3792 18340
rect 1780 18281 1808 18312
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 3620 18136 3648 18235
rect 3896 18213 3924 18380
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 5534 18408 5540 18420
rect 5316 18380 5540 18408
rect 5316 18368 5322 18380
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 5718 18368 5724 18420
rect 5776 18368 5782 18420
rect 10137 18411 10195 18417
rect 10137 18408 10149 18411
rect 6380 18380 10149 18408
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 6380 18340 6408 18380
rect 10137 18377 10149 18380
rect 10183 18377 10195 18411
rect 10137 18371 10195 18377
rect 10505 18411 10563 18417
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 14182 18408 14188 18420
rect 10551 18380 14188 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 15010 18368 15016 18420
rect 15068 18408 15074 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15068 18380 15669 18408
rect 15068 18368 15074 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 15749 18411 15807 18417
rect 15749 18377 15761 18411
rect 15795 18408 15807 18411
rect 17770 18408 17776 18420
rect 15795 18380 17776 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 18340 18380 18736 18408
rect 5675 18312 6408 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 6972 18312 7314 18340
rect 6972 18300 6978 18312
rect 8110 18300 8116 18352
rect 8168 18340 8174 18352
rect 9674 18340 9680 18352
rect 8168 18312 9680 18340
rect 8168 18300 8174 18312
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 11333 18343 11391 18349
rect 9784 18312 10916 18340
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9122 18272 9128 18284
rect 8803 18244 9128 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 9784 18272 9812 18312
rect 9456 18244 9812 18272
rect 10888 18272 10916 18312
rect 11333 18309 11345 18343
rect 11379 18340 11391 18343
rect 11790 18340 11796 18352
rect 11379 18312 11796 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 13909 18343 13967 18349
rect 13909 18309 13921 18343
rect 13955 18340 13967 18343
rect 13998 18340 14004 18352
rect 13955 18312 14004 18340
rect 13955 18309 13967 18312
rect 13909 18303 13967 18309
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 17313 18343 17371 18349
rect 17313 18309 17325 18343
rect 17359 18340 17371 18343
rect 18340 18340 18368 18380
rect 18708 18340 18736 18380
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19300 18380 19809 18408
rect 19300 18368 19306 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 22646 18408 22652 18420
rect 19797 18371 19855 18377
rect 20272 18380 22652 18408
rect 20070 18340 20076 18352
rect 17359 18312 18368 18340
rect 18432 18312 18644 18340
rect 18708 18312 20076 18340
rect 17359 18309 17371 18312
rect 17313 18303 17371 18309
rect 12069 18275 12127 18281
rect 12069 18272 12081 18275
rect 10888 18244 12081 18272
rect 9456 18232 9462 18244
rect 12069 18241 12081 18244
rect 12115 18272 12127 18275
rect 12526 18272 12532 18284
rect 12115 18244 12532 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 13078 18232 13084 18284
rect 13136 18232 13142 18284
rect 15856 18244 16068 18272
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 5905 18207 5963 18213
rect 5905 18204 5917 18207
rect 3881 18167 3939 18173
rect 3988 18176 5917 18204
rect 3988 18136 4016 18176
rect 5905 18173 5917 18176
rect 5951 18204 5963 18207
rect 5994 18204 6000 18216
rect 5951 18176 6000 18204
rect 5951 18173 5963 18176
rect 5905 18167 5963 18173
rect 5994 18164 6000 18176
rect 6052 18164 6058 18216
rect 6549 18207 6607 18213
rect 6549 18173 6561 18207
rect 6595 18173 6607 18207
rect 6549 18167 6607 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7282 18204 7288 18216
rect 6871 18176 7288 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 3620 18108 4016 18136
rect 4890 18096 4896 18148
rect 4948 18136 4954 18148
rect 6564 18136 6592 18167
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 9493 18207 9551 18213
rect 9493 18204 9505 18207
rect 7852 18176 9505 18204
rect 4948 18108 6592 18136
rect 4948 18096 4954 18108
rect 5258 18028 5264 18080
rect 5316 18028 5322 18080
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 5994 18068 6000 18080
rect 5684 18040 6000 18068
rect 5684 18028 5690 18040
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 6564 18068 6592 18108
rect 6914 18068 6920 18080
rect 6564 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18068 6978 18080
rect 7852 18068 7880 18176
rect 9493 18173 9505 18176
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 10594 18164 10600 18216
rect 10652 18164 10658 18216
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 8297 18139 8355 18145
rect 8297 18136 8309 18139
rect 7984 18108 8309 18136
rect 7984 18096 7990 18108
rect 8297 18105 8309 18108
rect 8343 18136 8355 18139
rect 8343 18108 8984 18136
rect 8343 18105 8355 18108
rect 8297 18099 8355 18105
rect 6972 18040 7880 18068
rect 8956 18068 8984 18108
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 9582 18136 9588 18148
rect 9088 18108 9588 18136
rect 9088 18096 9094 18108
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 10704 18068 10732 18167
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 12253 18207 12311 18213
rect 12253 18204 12265 18207
rect 11664 18176 12265 18204
rect 11664 18164 11670 18176
rect 12253 18173 12265 18176
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12986 18164 12992 18216
rect 13044 18204 13050 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 13044 18176 13185 18204
rect 13044 18164 13050 18176
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 12713 18139 12771 18145
rect 12713 18136 12725 18139
rect 10928 18108 12725 18136
rect 10928 18096 10934 18108
rect 12713 18105 12725 18108
rect 12759 18105 12771 18139
rect 12713 18099 12771 18105
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 13280 18136 13308 18167
rect 14550 18164 14556 18216
rect 14608 18204 14614 18216
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 14608 18176 14657 18204
rect 14608 18164 14614 18176
rect 14645 18173 14657 18176
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 14734 18164 14740 18216
rect 14792 18204 14798 18216
rect 15856 18204 15884 18244
rect 14792 18176 15884 18204
rect 14792 18164 14798 18176
rect 15930 18164 15936 18216
rect 15988 18164 15994 18216
rect 16040 18204 16068 18244
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 17092 18244 17233 18272
rect 17092 18232 17098 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 18432 18272 18460 18312
rect 17221 18235 17279 18241
rect 17420 18244 18460 18272
rect 18509 18275 18567 18281
rect 17420 18204 17448 18244
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18616 18272 18644 18312
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 19521 18275 19579 18281
rect 18616 18244 18736 18272
rect 18509 18235 18567 18241
rect 16040 18176 17448 18204
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 17497 18167 17555 18173
rect 12860 18108 13308 18136
rect 12860 18096 12866 18108
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 13504 18108 16528 18136
rect 13504 18096 13510 18108
rect 8956 18040 10732 18068
rect 6972 18028 6978 18040
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11609 18071 11667 18077
rect 11609 18068 11621 18071
rect 11480 18040 11621 18068
rect 11480 18028 11486 18040
rect 11609 18037 11621 18040
rect 11655 18068 11667 18071
rect 12434 18068 12440 18080
rect 11655 18040 12440 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14734 18068 14740 18080
rect 13872 18040 14740 18068
rect 13872 18028 13878 18040
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 15289 18071 15347 18077
rect 15289 18037 15301 18071
rect 15335 18068 15347 18071
rect 16114 18068 16120 18080
rect 15335 18040 16120 18068
rect 15335 18037 15347 18040
rect 15289 18031 15347 18037
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16356 18040 16405 18068
rect 16356 18028 16362 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16500 18068 16528 18108
rect 16850 18096 16856 18148
rect 16908 18096 16914 18148
rect 17512 18136 17540 18167
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18524 18204 18552 18235
rect 18288 18176 18552 18204
rect 18288 18164 18294 18176
rect 18598 18164 18604 18216
rect 18656 18164 18662 18216
rect 18708 18213 18736 18244
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 19978 18272 19984 18284
rect 19567 18244 19984 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 19978 18232 19984 18244
rect 20036 18272 20042 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20036 18244 20177 18272
rect 20036 18232 20042 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 19024 18176 19748 18204
rect 19024 18164 19030 18176
rect 19610 18136 19616 18148
rect 17512 18108 19616 18136
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 19720 18136 19748 18176
rect 19794 18164 19800 18216
rect 19852 18204 19858 18216
rect 20272 18213 20300 18380
rect 22646 18368 22652 18380
rect 22704 18368 22710 18420
rect 23198 18408 23204 18420
rect 23032 18380 23204 18408
rect 23032 18340 23060 18380
rect 23198 18368 23204 18380
rect 23256 18368 23262 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 25038 18408 25044 18420
rect 23440 18380 25044 18408
rect 23440 18368 23446 18380
rect 25038 18368 25044 18380
rect 25096 18408 25102 18420
rect 27157 18411 27215 18417
rect 25096 18380 25360 18408
rect 25096 18368 25102 18380
rect 23658 18340 23664 18352
rect 20824 18312 23060 18340
rect 23124 18312 23664 18340
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 19852 18176 20269 18204
rect 19852 18164 19858 18176
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 20346 18164 20352 18216
rect 20404 18164 20410 18216
rect 20824 18136 20852 18312
rect 23124 18281 23152 18312
rect 23658 18300 23664 18312
rect 23716 18300 23722 18352
rect 25332 18349 25360 18380
rect 27157 18377 27169 18411
rect 27203 18408 27215 18411
rect 27706 18408 27712 18420
rect 27203 18380 27712 18408
rect 27203 18377 27215 18380
rect 27157 18371 27215 18377
rect 27706 18368 27712 18380
rect 27764 18368 27770 18420
rect 29362 18408 29368 18420
rect 27816 18380 29368 18408
rect 25317 18343 25375 18349
rect 25317 18309 25329 18343
rect 25363 18309 25375 18343
rect 25317 18303 25375 18309
rect 25958 18300 25964 18352
rect 26016 18340 26022 18352
rect 27816 18340 27844 18380
rect 29362 18368 29368 18380
rect 29420 18368 29426 18420
rect 29822 18368 29828 18420
rect 29880 18368 29886 18420
rect 30745 18411 30803 18417
rect 30745 18377 30757 18411
rect 30791 18408 30803 18411
rect 37182 18408 37188 18420
rect 30791 18380 37188 18408
rect 30791 18377 30803 18380
rect 30745 18371 30803 18377
rect 37182 18368 37188 18380
rect 37240 18368 37246 18420
rect 28350 18340 28356 18352
rect 26016 18312 27844 18340
rect 28092 18312 28356 18340
rect 26016 18300 26022 18312
rect 28092 18284 28120 18312
rect 28350 18300 28356 18312
rect 28408 18300 28414 18352
rect 29638 18300 29644 18352
rect 29696 18340 29702 18352
rect 31573 18343 31631 18349
rect 31573 18340 31585 18343
rect 29696 18312 31585 18340
rect 29696 18300 29702 18312
rect 31573 18309 31585 18312
rect 31619 18340 31631 18343
rect 32125 18343 32183 18349
rect 32125 18340 32137 18343
rect 31619 18312 32137 18340
rect 31619 18309 31631 18312
rect 31573 18303 31631 18309
rect 32125 18309 32137 18312
rect 32171 18309 32183 18343
rect 32125 18303 32183 18309
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 21266 18164 21272 18216
rect 21324 18164 21330 18216
rect 19720 18108 20852 18136
rect 18141 18071 18199 18077
rect 18141 18068 18153 18071
rect 16500 18040 18153 18068
rect 16393 18031 16451 18037
rect 18141 18037 18153 18040
rect 18187 18037 18199 18071
rect 18141 18031 18199 18037
rect 19334 18028 19340 18080
rect 19392 18028 19398 18080
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 20346 18068 20352 18080
rect 19484 18040 20352 18068
rect 19484 18028 19490 18040
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20898 18068 20904 18080
rect 20496 18040 20904 18068
rect 20496 18028 20502 18040
rect 20898 18028 20904 18040
rect 20956 18028 20962 18080
rect 20993 18071 21051 18077
rect 20993 18037 21005 18071
rect 21039 18068 21051 18071
rect 21358 18068 21364 18080
rect 21039 18040 21364 18068
rect 21039 18037 21051 18040
rect 20993 18031 21051 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 22020 18068 22048 18235
rect 24394 18232 24400 18284
rect 24452 18272 24458 18284
rect 26786 18272 26792 18284
rect 24452 18244 26792 18272
rect 24452 18232 24458 18244
rect 26786 18232 26792 18244
rect 26844 18232 26850 18284
rect 28074 18232 28080 18284
rect 28132 18232 28138 18284
rect 29454 18232 29460 18284
rect 29512 18232 29518 18284
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18272 30711 18275
rect 31110 18272 31116 18284
rect 30699 18244 31116 18272
rect 30699 18241 30711 18244
rect 30653 18235 30711 18241
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 22649 18207 22707 18213
rect 22649 18173 22661 18207
rect 22695 18204 22707 18207
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 22695 18176 23397 18204
rect 22695 18173 22707 18176
rect 22649 18167 22707 18173
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 23750 18164 23756 18216
rect 23808 18204 23814 18216
rect 26053 18207 26111 18213
rect 26053 18204 26065 18207
rect 23808 18176 26065 18204
rect 23808 18164 23814 18176
rect 26053 18173 26065 18176
rect 26099 18173 26111 18207
rect 26053 18167 26111 18173
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18204 28411 18207
rect 30282 18204 30288 18216
rect 28399 18176 30288 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 30282 18164 30288 18176
rect 30340 18164 30346 18216
rect 30834 18164 30840 18216
rect 30892 18164 30898 18216
rect 24762 18096 24768 18148
rect 24820 18136 24826 18148
rect 24857 18139 24915 18145
rect 24857 18136 24869 18139
rect 24820 18108 24869 18136
rect 24820 18096 24826 18108
rect 24857 18105 24869 18108
rect 24903 18105 24915 18139
rect 24857 18099 24915 18105
rect 31754 18096 31760 18148
rect 31812 18096 31818 18148
rect 25314 18068 25320 18080
rect 22020 18040 25320 18068
rect 25314 18028 25320 18040
rect 25372 18068 25378 18080
rect 26510 18068 26516 18080
rect 25372 18040 26516 18068
rect 25372 18028 25378 18040
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 26697 18071 26755 18077
rect 26697 18037 26709 18071
rect 26743 18068 26755 18071
rect 26786 18068 26792 18080
rect 26743 18040 26792 18068
rect 26743 18037 26755 18040
rect 26697 18031 26755 18037
rect 26786 18028 26792 18040
rect 26844 18068 26850 18080
rect 27430 18068 27436 18080
rect 26844 18040 27436 18068
rect 26844 18028 26850 18040
rect 27430 18028 27436 18040
rect 27488 18068 27494 18080
rect 27709 18071 27767 18077
rect 27709 18068 27721 18071
rect 27488 18040 27721 18068
rect 27488 18028 27494 18040
rect 27709 18037 27721 18040
rect 27755 18068 27767 18071
rect 29454 18068 29460 18080
rect 27755 18040 29460 18068
rect 27755 18037 27767 18040
rect 27709 18031 27767 18037
rect 29454 18028 29460 18040
rect 29512 18028 29518 18080
rect 30282 18028 30288 18080
rect 30340 18028 30346 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 3418 17824 3424 17876
rect 3476 17824 3482 17876
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 10318 17864 10324 17876
rect 6236 17836 10324 17864
rect 6236 17824 6242 17836
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10502 17824 10508 17876
rect 10560 17824 10566 17876
rect 13814 17864 13820 17876
rect 11072 17836 13820 17864
rect 6730 17796 6736 17808
rect 2746 17768 6736 17796
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 2746 17660 2774 17768
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 8757 17799 8815 17805
rect 6840 17768 8340 17796
rect 3878 17688 3884 17740
rect 3936 17728 3942 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 3936 17700 4445 17728
rect 3936 17688 3942 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4614 17688 4620 17740
rect 4672 17728 4678 17740
rect 6273 17731 6331 17737
rect 6273 17728 6285 17731
rect 4672 17700 6285 17728
rect 4672 17688 4678 17700
rect 6273 17697 6285 17700
rect 6319 17697 6331 17731
rect 6273 17691 6331 17697
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6840 17728 6868 17768
rect 6604 17700 6868 17728
rect 6604 17688 6610 17700
rect 8110 17688 8116 17740
rect 8168 17728 8174 17740
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 8168 17700 8217 17728
rect 8168 17688 8174 17700
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8312 17728 8340 17768
rect 8757 17765 8769 17799
rect 8803 17796 8815 17799
rect 10520 17796 10548 17824
rect 8803 17768 10548 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 11072 17737 11100 17836
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 13909 17867 13967 17873
rect 13909 17833 13921 17867
rect 13955 17833 13967 17867
rect 13909 17827 13967 17833
rect 13924 17796 13952 17827
rect 14458 17824 14464 17876
rect 14516 17824 14522 17876
rect 14826 17824 14832 17876
rect 14884 17824 14890 17876
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 15896 17836 18061 17864
rect 15896 17824 15902 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 18049 17827 18107 17833
rect 13998 17796 14004 17808
rect 13924 17768 14004 17796
rect 13998 17756 14004 17768
rect 14056 17796 14062 17808
rect 15194 17796 15200 17808
rect 14056 17768 15200 17796
rect 14056 17756 14062 17768
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 18064 17796 18092 17827
rect 19242 17824 19248 17876
rect 19300 17864 19306 17876
rect 19300 17836 21404 17864
rect 19300 17824 19306 17836
rect 20438 17796 20444 17808
rect 18064 17768 20444 17796
rect 20438 17756 20444 17768
rect 20496 17756 20502 17808
rect 20898 17756 20904 17808
rect 20956 17796 20962 17808
rect 20956 17768 21312 17796
rect 20956 17756 20962 17768
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 8312 17700 10977 17728
rect 8205 17691 8263 17697
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 11057 17731 11115 17737
rect 11057 17697 11069 17731
rect 11103 17697 11115 17731
rect 11057 17691 11115 17697
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 11606 17728 11612 17740
rect 11388 17700 11612 17728
rect 11388 17688 11394 17700
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 14550 17728 14556 17740
rect 11756 17700 14556 17728
rect 11756 17688 11762 17700
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 16264 17700 16313 17728
rect 16264 17688 16270 17700
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 20622 17728 20628 17740
rect 16623 17700 20628 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 21284 17737 21312 17768
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20864 17700 21189 17728
rect 20864 17688 20870 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17697 21327 17731
rect 21376 17728 21404 17836
rect 21726 17824 21732 17876
rect 21784 17824 21790 17876
rect 21910 17824 21916 17876
rect 21968 17824 21974 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 24084 17836 24685 17864
rect 24084 17824 24090 17836
rect 24673 17833 24685 17836
rect 24719 17864 24731 17867
rect 24762 17864 24768 17876
rect 24719 17836 24768 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 26510 17824 26516 17876
rect 26568 17864 26574 17876
rect 26697 17867 26755 17873
rect 26697 17864 26709 17867
rect 26568 17836 26709 17864
rect 26568 17824 26574 17836
rect 26697 17833 26709 17836
rect 26743 17833 26755 17867
rect 26697 17827 26755 17833
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 27672 17836 28764 17864
rect 27672 17824 27678 17836
rect 28736 17740 28764 17836
rect 28902 17824 28908 17876
rect 28960 17864 28966 17876
rect 30834 17864 30840 17876
rect 28960 17836 30840 17864
rect 28960 17824 28966 17836
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 31110 17824 31116 17876
rect 31168 17864 31174 17876
rect 31297 17867 31355 17873
rect 31297 17864 31309 17867
rect 31168 17836 31309 17864
rect 31168 17824 31174 17836
rect 31297 17833 31309 17836
rect 31343 17833 31355 17867
rect 31297 17827 31355 17833
rect 30374 17756 30380 17808
rect 30432 17796 30438 17808
rect 32490 17796 32496 17808
rect 30432 17768 32496 17796
rect 30432 17756 30438 17768
rect 32490 17756 32496 17768
rect 32548 17756 32554 17808
rect 23750 17728 23756 17740
rect 21376 17700 23756 17728
rect 21269 17691 21327 17697
rect 23750 17688 23756 17700
rect 23808 17728 23814 17740
rect 24397 17731 24455 17737
rect 24397 17728 24409 17731
rect 23808 17700 24409 17728
rect 23808 17688 23814 17700
rect 24397 17697 24409 17700
rect 24443 17697 24455 17731
rect 24397 17691 24455 17697
rect 1811 17632 2774 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 4062 17620 4068 17672
rect 4120 17620 4126 17672
rect 5997 17663 6055 17669
rect 5997 17629 6009 17663
rect 6043 17660 6055 17663
rect 7006 17660 7012 17672
rect 6043 17632 7012 17660
rect 6043 17629 6055 17632
rect 5997 17623 6055 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17660 8079 17663
rect 8067 17632 11100 17660
rect 8067 17629 8079 17632
rect 8021 17623 8079 17629
rect 1394 17552 1400 17604
rect 1452 17592 1458 17604
rect 4798 17592 4804 17604
rect 1452 17564 4804 17592
rect 1452 17552 1458 17564
rect 4798 17552 4804 17564
rect 4856 17592 4862 17604
rect 6638 17592 6644 17604
rect 4856 17564 6644 17592
rect 4856 17552 4862 17564
rect 6638 17552 6644 17564
rect 6696 17552 6702 17604
rect 6822 17552 6828 17604
rect 6880 17592 6886 17604
rect 6880 17564 9076 17592
rect 6880 17552 6886 17564
rect 3605 17527 3663 17533
rect 3605 17493 3617 17527
rect 3651 17524 3663 17527
rect 3878 17524 3884 17536
rect 3651 17496 3884 17524
rect 3651 17493 3663 17496
rect 3605 17487 3663 17493
rect 3878 17484 3884 17496
rect 3936 17524 3942 17536
rect 6546 17524 6552 17536
rect 3936 17496 6552 17524
rect 3936 17484 3942 17496
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 7156 17496 7665 17524
rect 7156 17484 7162 17496
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 7653 17487 7711 17493
rect 8113 17527 8171 17533
rect 8113 17493 8125 17527
rect 8159 17524 8171 17527
rect 8202 17524 8208 17536
rect 8159 17496 8208 17524
rect 8159 17493 8171 17496
rect 8113 17487 8171 17493
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 9048 17524 9076 17564
rect 9122 17552 9128 17604
rect 9180 17552 9186 17604
rect 9858 17552 9864 17604
rect 9916 17552 9922 17604
rect 10413 17595 10471 17601
rect 10413 17561 10425 17595
rect 10459 17592 10471 17595
rect 10459 17564 10824 17592
rect 10459 17561 10471 17564
rect 10413 17555 10471 17561
rect 10796 17536 10824 17564
rect 9674 17524 9680 17536
rect 9048 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 10594 17524 10600 17536
rect 10551 17496 10600 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10836 17496 10885 17524
rect 10836 17484 10842 17496
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 11072 17524 11100 17632
rect 13630 17620 13636 17672
rect 13688 17660 13694 17672
rect 15197 17663 15255 17669
rect 15197 17660 15209 17663
rect 13688 17632 15209 17660
rect 13688 17620 13694 17632
rect 15197 17629 15209 17632
rect 15243 17660 15255 17663
rect 15838 17660 15844 17672
rect 15243 17632 15844 17660
rect 15243 17629 15255 17632
rect 15197 17623 15255 17629
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17660 19395 17663
rect 19426 17660 19432 17672
rect 19383 17632 19432 17660
rect 19383 17629 19395 17632
rect 19337 17623 19395 17629
rect 19426 17620 19432 17632
rect 19484 17620 19490 17672
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20128 17632 20760 17660
rect 20128 17620 20134 17632
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 11977 17595 12035 17601
rect 11977 17592 11989 17595
rect 11388 17564 11989 17592
rect 11388 17552 11394 17564
rect 11977 17561 11989 17564
rect 12023 17561 12035 17595
rect 11977 17555 12035 17561
rect 12434 17552 12440 17604
rect 12492 17552 12498 17604
rect 13814 17592 13820 17604
rect 13372 17564 13820 17592
rect 13372 17524 13400 17564
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 13906 17552 13912 17604
rect 13964 17592 13970 17604
rect 14369 17595 14427 17601
rect 14369 17592 14381 17595
rect 13964 17564 14381 17592
rect 13964 17552 13970 17564
rect 14369 17561 14381 17564
rect 14415 17561 14427 17595
rect 14369 17555 14427 17561
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 18601 17595 18659 17601
rect 16540 17564 17066 17592
rect 16540 17552 16546 17564
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 20162 17592 20168 17604
rect 18647 17564 20168 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 20162 17552 20168 17564
rect 20220 17552 20226 17604
rect 20254 17552 20260 17604
rect 20312 17552 20318 17604
rect 11072 17496 13400 17524
rect 13449 17527 13507 17533
rect 10873 17487 10931 17493
rect 13449 17493 13461 17527
rect 13495 17524 13507 17527
rect 14090 17524 14096 17536
rect 13495 17496 14096 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14458 17524 14464 17536
rect 14332 17496 14464 17524
rect 14332 17484 14338 17496
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 15838 17484 15844 17536
rect 15896 17484 15902 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 20732 17533 20760 17632
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 21140 17632 22293 17660
rect 21140 17620 21146 17632
rect 22281 17629 22293 17632
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 21692 17564 22569 17592
rect 21692 17552 21698 17564
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 23842 17592 23848 17604
rect 23782 17564 23848 17592
rect 22557 17555 22615 17561
rect 23842 17552 23848 17564
rect 23900 17592 23906 17604
rect 24302 17592 24308 17604
rect 23900 17564 24308 17592
rect 23900 17552 23906 17564
rect 24302 17552 24308 17564
rect 24360 17552 24366 17604
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 17276 17496 18705 17524
rect 17276 17484 17282 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17493 20775 17527
rect 20717 17487 20775 17493
rect 21085 17527 21143 17533
rect 21085 17493 21097 17527
rect 21131 17524 21143 17527
rect 21358 17524 21364 17536
rect 21131 17496 21364 17524
rect 21131 17493 21143 17496
rect 21085 17487 21143 17493
rect 21358 17484 21364 17496
rect 21416 17524 21422 17536
rect 21818 17524 21824 17536
rect 21416 17496 21824 17524
rect 21416 17484 21422 17496
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 21910 17484 21916 17536
rect 21968 17524 21974 17536
rect 22462 17524 22468 17536
rect 21968 17496 22468 17524
rect 21968 17484 21974 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 24029 17527 24087 17533
rect 24029 17524 24041 17527
rect 23348 17496 24041 17524
rect 23348 17484 23354 17496
rect 24029 17493 24041 17496
rect 24075 17524 24087 17527
rect 24118 17524 24124 17536
rect 24075 17496 24124 17524
rect 24075 17493 24087 17496
rect 24029 17487 24087 17493
rect 24118 17484 24124 17496
rect 24176 17484 24182 17536
rect 24412 17524 24440 17691
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 27157 17731 27215 17737
rect 27157 17728 27169 17731
rect 25004 17700 27169 17728
rect 25004 17688 25010 17700
rect 27157 17697 27169 17700
rect 27203 17728 27215 17731
rect 27798 17728 27804 17740
rect 27203 17700 27804 17728
rect 27203 17697 27215 17700
rect 27157 17691 27215 17697
rect 27798 17688 27804 17700
rect 27856 17728 27862 17740
rect 28074 17728 28080 17740
rect 27856 17700 28080 17728
rect 27856 17688 27862 17700
rect 28074 17688 28080 17700
rect 28132 17688 28138 17740
rect 28718 17688 28724 17740
rect 28776 17728 28782 17740
rect 28776 17700 29592 17728
rect 28776 17688 28782 17700
rect 29273 17663 29331 17669
rect 29273 17660 29285 17663
rect 28566 17632 29285 17660
rect 29273 17629 29285 17632
rect 29319 17660 29331 17663
rect 29454 17660 29460 17672
rect 29319 17632 29460 17660
rect 29319 17629 29331 17632
rect 29273 17623 29331 17629
rect 29454 17620 29460 17632
rect 29512 17620 29518 17672
rect 29564 17660 29592 17700
rect 30006 17688 30012 17740
rect 30064 17728 30070 17740
rect 30285 17731 30343 17737
rect 30285 17728 30297 17731
rect 30064 17700 30297 17728
rect 30064 17688 30070 17700
rect 30285 17697 30297 17700
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 30837 17731 30895 17737
rect 30837 17697 30849 17731
rect 30883 17728 30895 17731
rect 31294 17728 31300 17740
rect 30883 17700 31300 17728
rect 30883 17697 30895 17700
rect 30837 17691 30895 17697
rect 31294 17688 31300 17700
rect 31352 17688 31358 17740
rect 31018 17660 31024 17672
rect 29564 17632 31024 17660
rect 31018 17620 31024 17632
rect 31076 17620 31082 17672
rect 31128 17632 41414 17660
rect 24854 17552 24860 17604
rect 24912 17592 24918 17604
rect 25225 17595 25283 17601
rect 25225 17592 25237 17595
rect 24912 17564 25237 17592
rect 24912 17552 24918 17564
rect 25225 17561 25237 17564
rect 25271 17561 25283 17595
rect 26786 17592 26792 17604
rect 26450 17564 26792 17592
rect 25225 17555 25283 17561
rect 26786 17552 26792 17564
rect 26844 17552 26850 17604
rect 27433 17595 27491 17601
rect 27433 17561 27445 17595
rect 27479 17592 27491 17595
rect 27706 17592 27712 17604
rect 27479 17564 27712 17592
rect 27479 17561 27491 17564
rect 27433 17555 27491 17561
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 31128 17601 31156 17632
rect 30101 17595 30159 17601
rect 30101 17592 30113 17595
rect 28736 17564 30113 17592
rect 28736 17524 28764 17564
rect 30101 17561 30113 17564
rect 30147 17592 30159 17595
rect 31113 17595 31171 17601
rect 31113 17592 31125 17595
rect 30147 17564 31125 17592
rect 30147 17561 30159 17564
rect 30101 17555 30159 17561
rect 31113 17561 31125 17564
rect 31159 17561 31171 17595
rect 41386 17592 41414 17632
rect 45462 17592 45468 17604
rect 41386 17564 45468 17592
rect 31113 17555 31171 17561
rect 45462 17552 45468 17564
rect 45520 17552 45526 17604
rect 24412 17496 28764 17524
rect 29362 17484 29368 17536
rect 29420 17524 29426 17536
rect 29733 17527 29791 17533
rect 29733 17524 29745 17527
rect 29420 17496 29745 17524
rect 29420 17484 29426 17496
rect 29733 17493 29745 17496
rect 29779 17493 29791 17527
rect 29733 17487 29791 17493
rect 30190 17484 30196 17536
rect 30248 17524 30254 17536
rect 30929 17527 30987 17533
rect 30929 17524 30941 17527
rect 30248 17496 30941 17524
rect 30248 17484 30254 17496
rect 30929 17493 30941 17496
rect 30975 17524 30987 17527
rect 47026 17524 47032 17536
rect 30975 17496 47032 17524
rect 30975 17493 30987 17496
rect 30929 17487 30987 17493
rect 47026 17484 47032 17496
rect 47084 17484 47090 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 7193 17323 7251 17329
rect 7193 17320 7205 17323
rect 5592 17292 7205 17320
rect 5592 17280 5598 17292
rect 7193 17289 7205 17292
rect 7239 17289 7251 17323
rect 7193 17283 7251 17289
rect 7285 17323 7343 17329
rect 7285 17289 7297 17323
rect 7331 17320 7343 17323
rect 9214 17320 9220 17332
rect 7331 17292 9220 17320
rect 7331 17289 7343 17292
rect 7285 17283 7343 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9456 17292 9597 17320
rect 9456 17280 9462 17292
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 9585 17283 9643 17289
rect 9674 17280 9680 17332
rect 9732 17280 9738 17332
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 20254 17320 20260 17332
rect 10376 17292 12434 17320
rect 10376 17280 10382 17292
rect 4246 17212 4252 17264
rect 4304 17252 4310 17264
rect 4341 17255 4399 17261
rect 4341 17252 4353 17255
rect 4304 17224 4353 17252
rect 4304 17212 4310 17224
rect 4341 17221 4353 17224
rect 4387 17221 4399 17255
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 4341 17215 4399 17221
rect 5552 17224 11989 17252
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 5552 17184 5580 17224
rect 11977 17221 11989 17224
rect 12023 17221 12035 17255
rect 12406 17252 12434 17292
rect 13740 17292 20260 17320
rect 13354 17252 13360 17264
rect 12406 17224 13360 17252
rect 11977 17215 12035 17221
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 13740 17261 13768 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 22557 17323 22615 17329
rect 22557 17320 22569 17323
rect 21324 17292 22569 17320
rect 21324 17280 21330 17292
rect 22557 17289 22569 17292
rect 22603 17289 22615 17323
rect 22557 17283 22615 17289
rect 22649 17323 22707 17329
rect 22649 17289 22661 17323
rect 22695 17320 22707 17323
rect 30282 17320 30288 17332
rect 22695 17292 30288 17320
rect 22695 17289 22707 17292
rect 22649 17283 22707 17289
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 13725 17255 13783 17261
rect 13725 17221 13737 17255
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 15562 17252 15568 17264
rect 14240 17224 15568 17252
rect 14240 17212 14246 17224
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 15838 17212 15844 17264
rect 15896 17252 15902 17264
rect 18417 17255 18475 17261
rect 18417 17252 18429 17255
rect 15896 17224 18429 17252
rect 15896 17212 15902 17224
rect 18417 17221 18429 17224
rect 18463 17221 18475 17255
rect 18417 17215 18475 17221
rect 21818 17212 21824 17264
rect 21876 17212 21882 17264
rect 23293 17255 23351 17261
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 23474 17252 23480 17264
rect 23339 17224 23480 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 23474 17212 23480 17224
rect 23532 17252 23538 17264
rect 23934 17252 23940 17264
rect 23532 17224 23940 17252
rect 23532 17212 23538 17224
rect 23934 17212 23940 17224
rect 23992 17212 23998 17264
rect 24026 17212 24032 17264
rect 24084 17212 24090 17264
rect 24946 17252 24952 17264
rect 24780 17224 24952 17252
rect 3651 17156 5580 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5736 17156 6592 17184
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 5736 17125 5764 17156
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 2924 17088 5733 17116
rect 2924 17076 2930 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 6564 17116 6592 17156
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6696 17156 7512 17184
rect 6696 17144 6702 17156
rect 7377 17119 7435 17125
rect 6564 17088 7052 17116
rect 5813 17079 5871 17085
rect 4890 17008 4896 17060
rect 4948 17048 4954 17060
rect 5828 17048 5856 17079
rect 4948 17020 5856 17048
rect 4948 17008 4954 17020
rect 6362 17008 6368 17060
rect 6420 17048 6426 17060
rect 6825 17051 6883 17057
rect 6825 17048 6837 17051
rect 6420 17020 6837 17048
rect 6420 17008 6426 17020
rect 6825 17017 6837 17020
rect 6871 17017 6883 17051
rect 6825 17011 6883 17017
rect 5261 16983 5319 16989
rect 5261 16949 5273 16983
rect 5307 16980 5319 16983
rect 5534 16980 5540 16992
rect 5307 16952 5540 16980
rect 5307 16949 5319 16952
rect 5261 16943 5319 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 6178 16940 6184 16992
rect 6236 16980 6242 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6236 16952 6469 16980
rect 6236 16940 6242 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 7024 16980 7052 17088
rect 7377 17085 7389 17119
rect 7423 17085 7435 17119
rect 7484 17116 7512 17156
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 9950 17184 9956 17196
rect 8588 17156 9956 17184
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 7484 17088 8493 17116
rect 7377 17079 7435 17085
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 7282 17008 7288 17060
rect 7340 17048 7346 17060
rect 7392 17048 7420 17079
rect 8588 17048 8616 17156
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 10827 17156 11376 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17085 8723 17119
rect 8665 17079 8723 17085
rect 7340 17020 8616 17048
rect 8680 17048 8708 17079
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9030 17116 9036 17128
rect 8904 17088 9036 17116
rect 8904 17076 8910 17088
rect 9030 17076 9036 17088
rect 9088 17116 9094 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9088 17088 9781 17116
rect 9088 17076 9094 17088
rect 9769 17085 9781 17088
rect 9815 17116 9827 17119
rect 10226 17116 10232 17128
rect 9815 17088 10232 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10376 17088 10885 17116
rect 10376 17076 10382 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 8680 17020 9812 17048
rect 7340 17008 7346 17020
rect 9784 16992 9812 17020
rect 10686 17008 10692 17060
rect 10744 17048 10750 17060
rect 10980 17048 11008 17079
rect 10744 17020 11008 17048
rect 10744 17008 10750 17020
rect 7926 16980 7932 16992
rect 7024 16952 7932 16980
rect 6457 16943 6515 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 8021 16983 8079 16989
rect 8021 16949 8033 16983
rect 8067 16980 8079 16983
rect 8202 16980 8208 16992
rect 8067 16952 8208 16980
rect 8067 16949 8079 16952
rect 8021 16943 8079 16949
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 8352 16952 9229 16980
rect 8352 16940 8358 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 10870 16940 10876 16992
rect 10928 16980 10934 16992
rect 11072 16980 11100 17156
rect 11348 17116 11376 17156
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11480 17156 11805 17184
rect 11480 17144 11486 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12124 17156 12817 17184
rect 12124 17144 12130 17156
rect 12805 17153 12817 17156
rect 12851 17153 12863 17187
rect 14090 17184 14096 17196
rect 12805 17147 12863 17153
rect 13004 17156 14096 17184
rect 12618 17116 12624 17128
rect 11348 17088 12624 17116
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 12894 17076 12900 17128
rect 12952 17076 12958 17128
rect 13004 17125 13032 17156
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14332 17156 14749 17184
rect 14332 17144 14338 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14826 17144 14832 17196
rect 14884 17144 14890 17196
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 16724 17156 17233 17184
rect 16724 17144 16730 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19550 17156 20177 17184
rect 17221 17147 17279 17153
rect 20165 17153 20177 17156
rect 20211 17184 20223 17187
rect 20530 17184 20536 17196
rect 20211 17156 20536 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 24780 17193 24808 17224
rect 24946 17212 24952 17224
rect 25004 17212 25010 17264
rect 26786 17252 26792 17264
rect 26266 17224 26792 17252
rect 26786 17212 26792 17224
rect 26844 17212 26850 17264
rect 29454 17252 29460 17264
rect 29394 17224 29460 17252
rect 29454 17212 29460 17224
rect 29512 17252 29518 17264
rect 30009 17255 30067 17261
rect 30009 17252 30021 17255
rect 29512 17224 30021 17252
rect 29512 17212 29518 17224
rect 30009 17221 30021 17224
rect 30055 17252 30067 17255
rect 31294 17252 31300 17264
rect 30055 17224 31300 17252
rect 30055 17221 30067 17224
rect 30009 17215 30067 17221
rect 31294 17212 31300 17224
rect 31352 17212 31358 17264
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 24765 17187 24823 17193
rect 20809 17147 20867 17153
rect 22572 17156 22876 17184
rect 12989 17119 13047 17125
rect 12989 17085 13001 17119
rect 13035 17085 13047 17119
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 12989 17079 13047 17085
rect 13096 17088 14933 17116
rect 12434 17008 12440 17060
rect 12492 17008 12498 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 13096 17048 13124 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 17313 17119 17371 17125
rect 17313 17116 17325 17119
rect 15988 17088 17325 17116
rect 15988 17076 15994 17088
rect 17313 17085 17325 17088
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17116 17555 17119
rect 17770 17116 17776 17128
rect 17543 17088 17776 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 12584 17020 13124 17048
rect 12584 17008 12590 17020
rect 13722 17008 13728 17060
rect 13780 17048 13786 17060
rect 16758 17048 16764 17060
rect 13780 17020 16764 17048
rect 13780 17008 13786 17020
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 18156 17048 18184 17079
rect 19610 17076 19616 17128
rect 19668 17116 19674 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19668 17088 19901 17116
rect 19668 17076 19674 17088
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 20824 17116 20852 17147
rect 22572 17116 22600 17156
rect 22848 17125 22876 17156
rect 24765 17153 24777 17187
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 27798 17144 27804 17196
rect 27856 17184 27862 17196
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27856 17156 27905 17184
rect 27856 17144 27862 17156
rect 27893 17153 27905 17156
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 20824 17088 22600 17116
rect 22833 17119 22891 17125
rect 19889 17079 19947 17085
rect 22833 17085 22845 17119
rect 22879 17116 22891 17119
rect 22879 17088 23796 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 17184 17020 18184 17048
rect 17184 17008 17190 17020
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 19852 17020 21036 17048
rect 19852 17008 19858 17020
rect 10928 16952 11100 16980
rect 10928 16940 10934 16952
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 13446 16980 13452 16992
rect 11848 16952 13452 16980
rect 11848 16940 11854 16952
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 13814 16940 13820 16992
rect 13872 16940 13878 16992
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14056 16952 14381 16980
rect 14056 16940 14062 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 14369 16943 14427 16949
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15436 16952 16313 16980
rect 15436 16940 15442 16952
rect 16301 16949 16313 16952
rect 16347 16949 16359 16983
rect 16301 16943 16359 16949
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16632 16952 16865 16980
rect 16632 16940 16638 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 20070 16980 20076 16992
rect 17092 16952 20076 16980
rect 17092 16940 17098 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20898 16980 20904 16992
rect 20680 16952 20904 16980
rect 20680 16940 20686 16952
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21008 16980 21036 17020
rect 21174 17008 21180 17060
rect 21232 17048 21238 17060
rect 22189 17051 22247 17057
rect 22189 17048 22201 17051
rect 21232 17020 22201 17048
rect 21232 17008 21238 17020
rect 22189 17017 22201 17020
rect 22235 17017 22247 17051
rect 22189 17011 22247 17017
rect 21453 16983 21511 16989
rect 21453 16980 21465 16983
rect 21008 16952 21465 16980
rect 21453 16949 21465 16952
rect 21499 16949 21511 16983
rect 21453 16943 21511 16949
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 21910 16980 21916 16992
rect 21784 16952 21916 16980
rect 21784 16940 21790 16952
rect 21910 16940 21916 16952
rect 21968 16980 21974 16992
rect 23474 16980 23480 16992
rect 21968 16952 23480 16980
rect 21968 16940 21974 16952
rect 23474 16940 23480 16952
rect 23532 16940 23538 16992
rect 23566 16940 23572 16992
rect 23624 16940 23630 16992
rect 23768 16980 23796 17088
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23992 17088 24133 17116
rect 23992 17076 23998 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24121 17079 24179 17085
rect 25041 17119 25099 17125
rect 25041 17085 25053 17119
rect 25087 17116 25099 17119
rect 25087 17088 26188 17116
rect 25087 17085 25099 17088
rect 25041 17079 25099 17085
rect 26160 17060 26188 17088
rect 27246 17076 27252 17128
rect 27304 17076 27310 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 30006 17116 30012 17128
rect 28215 17088 30012 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 30006 17076 30012 17088
rect 30064 17076 30070 17128
rect 26142 17008 26148 17060
rect 26200 17008 26206 17060
rect 32858 17008 32864 17060
rect 32916 17048 32922 17060
rect 34514 17048 34520 17060
rect 32916 17020 34520 17048
rect 32916 17008 32922 17020
rect 34514 17008 34520 17020
rect 34572 17008 34578 17060
rect 26513 16983 26571 16989
rect 26513 16980 26525 16983
rect 23768 16952 26525 16980
rect 26513 16949 26525 16952
rect 26559 16949 26571 16983
rect 26513 16943 26571 16949
rect 27522 16940 27528 16992
rect 27580 16980 27586 16992
rect 29641 16983 29699 16989
rect 29641 16980 29653 16983
rect 27580 16952 29653 16980
rect 27580 16940 27586 16952
rect 29641 16949 29653 16952
rect 29687 16949 29699 16983
rect 29641 16943 29699 16949
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 3418 16736 3424 16788
rect 3476 16736 3482 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 6086 16776 6092 16788
rect 5132 16748 6092 16776
rect 5132 16736 5138 16748
rect 6086 16736 6092 16748
rect 6144 16776 6150 16788
rect 6144 16748 8248 16776
rect 6144 16736 6150 16748
rect 3513 16711 3571 16717
rect 3513 16708 3525 16711
rect 2746 16680 3525 16708
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 2746 16640 2774 16680
rect 3513 16677 3525 16680
rect 3559 16708 3571 16711
rect 8220 16708 8248 16748
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 10321 16779 10379 16785
rect 10321 16776 10333 16779
rect 9732 16748 10333 16776
rect 9732 16736 9738 16748
rect 10321 16745 10333 16748
rect 10367 16776 10379 16779
rect 12066 16776 12072 16788
rect 10367 16748 12072 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 14182 16776 14188 16788
rect 12308 16748 14188 16776
rect 12308 16736 12314 16748
rect 3559 16680 8064 16708
rect 8220 16680 8432 16708
rect 3559 16677 3571 16680
rect 3513 16671 3571 16677
rect 2280 16612 2774 16640
rect 2280 16600 2286 16612
rect 3326 16600 3332 16652
rect 3384 16640 3390 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 3384 16612 6193 16640
rect 3384 16600 3390 16612
rect 6181 16609 6193 16612
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 7098 16600 7104 16652
rect 7156 16600 7162 16652
rect 7282 16600 7288 16652
rect 7340 16600 7346 16652
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 4065 16575 4123 16581
rect 1811 16544 2774 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 2501 16467 2559 16473
rect 2746 16436 2774 16544
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 4080 16504 4108 16535
rect 4706 16532 4712 16584
rect 4764 16572 4770 16584
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4764 16544 4905 16572
rect 4764 16532 4770 16544
rect 4893 16541 4905 16544
rect 4939 16541 4951 16575
rect 7834 16572 7840 16584
rect 4893 16535 4951 16541
rect 5000 16544 7840 16572
rect 5000 16504 5028 16544
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 8036 16572 8064 16680
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8404 16649 8432 16680
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 9398 16708 9404 16720
rect 8720 16680 9404 16708
rect 8720 16668 8726 16680
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 11793 16711 11851 16717
rect 9600 16680 10272 16708
rect 9600 16649 9628 16680
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8168 16612 8309 16640
rect 8168 16600 8174 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16609 8447 16643
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 8389 16603 8447 16609
rect 8496 16612 9597 16640
rect 8496 16572 8524 16612
rect 9585 16609 9597 16612
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9766 16600 9772 16652
rect 9824 16600 9830 16652
rect 10244 16649 10272 16680
rect 11793 16677 11805 16711
rect 11839 16708 11851 16711
rect 11839 16680 12388 16708
rect 11839 16677 11851 16680
rect 11793 16671 11851 16677
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 10275 16612 12265 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 8036 16544 8524 16572
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 9493 16575 9551 16581
rect 9493 16572 9505 16575
rect 8812 16544 9505 16572
rect 8812 16532 8818 16544
rect 9493 16541 9505 16544
rect 9539 16541 9551 16575
rect 9784 16572 9812 16600
rect 10594 16572 10600 16584
rect 9784 16544 10600 16572
rect 9493 16535 9551 16541
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 11790 16572 11796 16584
rect 10735 16544 11796 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 12161 16575 12219 16581
rect 12161 16572 12173 16575
rect 12124 16544 12173 16572
rect 12124 16532 12130 16544
rect 12161 16541 12173 16544
rect 12207 16541 12219 16575
rect 12360 16572 12388 16680
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12544 16640 12572 16748
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14458 16736 14464 16788
rect 14516 16736 14522 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 14700 16748 16313 16776
rect 14700 16736 14706 16748
rect 16301 16745 16313 16748
rect 16347 16776 16359 16779
rect 18966 16776 18972 16788
rect 16347 16748 18972 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 23014 16776 23020 16788
rect 20128 16748 23020 16776
rect 20128 16736 20134 16748
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23290 16736 23296 16788
rect 23348 16736 23354 16788
rect 24118 16736 24124 16788
rect 24176 16776 24182 16788
rect 24176 16748 29868 16776
rect 24176 16736 24182 16748
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 16942 16708 16948 16720
rect 13035 16680 16948 16708
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 18506 16668 18512 16720
rect 18564 16708 18570 16720
rect 18785 16711 18843 16717
rect 18785 16708 18797 16711
rect 18564 16680 18797 16708
rect 18564 16668 18570 16680
rect 18785 16677 18797 16680
rect 18831 16708 18843 16711
rect 18874 16708 18880 16720
rect 18831 16680 18880 16708
rect 18831 16677 18843 16680
rect 18785 16671 18843 16677
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 29730 16708 29736 16720
rect 20772 16680 26280 16708
rect 20772 16668 20778 16680
rect 12483 16612 12572 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 13262 16640 13268 16652
rect 12676 16612 13268 16640
rect 12676 16600 12682 16612
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13446 16600 13452 16652
rect 13504 16600 13510 16652
rect 13630 16600 13636 16652
rect 13688 16600 13694 16652
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 14424 16612 15608 16640
rect 14424 16600 14430 16612
rect 15010 16572 15016 16584
rect 12360 16544 15016 16572
rect 12161 16535 12219 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 15580 16572 15608 16612
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 16298 16640 16304 16652
rect 15712 16612 16304 16640
rect 15712 16600 15718 16612
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16408 16612 18552 16640
rect 16117 16575 16175 16581
rect 15580 16544 16068 16572
rect 4080 16476 5028 16504
rect 5997 16507 6055 16513
rect 5997 16473 6009 16507
rect 6043 16504 6055 16507
rect 6270 16504 6276 16516
rect 6043 16476 6276 16504
rect 6043 16473 6055 16476
rect 5997 16467 6055 16473
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7156 16476 8217 16504
rect 7156 16464 7162 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 8570 16464 8576 16516
rect 8628 16504 8634 16516
rect 9858 16504 9864 16516
rect 8628 16476 9864 16504
rect 8628 16464 8634 16476
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 11422 16504 11428 16516
rect 10192 16476 11428 16504
rect 10192 16464 10198 16476
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 13538 16504 13544 16516
rect 12492 16476 13544 16504
rect 12492 16464 12498 16476
rect 13538 16464 13544 16476
rect 13596 16464 13602 16516
rect 14369 16507 14427 16513
rect 14369 16473 14381 16507
rect 14415 16504 14427 16507
rect 14642 16504 14648 16516
rect 14415 16476 14648 16504
rect 14415 16473 14427 16476
rect 14369 16467 14427 16473
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 15381 16507 15439 16513
rect 15381 16473 15393 16507
rect 15427 16504 15439 16507
rect 15746 16504 15752 16516
rect 15427 16476 15752 16504
rect 15427 16473 15439 16476
rect 15381 16467 15439 16473
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 16040 16504 16068 16544
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16206 16572 16212 16584
rect 16163 16544 16212 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16408 16504 16436 16612
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16572 16727 16575
rect 16758 16572 16764 16584
rect 16715 16544 16764 16572
rect 16715 16541 16727 16544
rect 16669 16535 16727 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 18524 16572 18552 16612
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18656 16612 19073 16640
rect 18656 16600 18662 16612
rect 19061 16609 19073 16612
rect 19107 16640 19119 16643
rect 19150 16640 19156 16652
rect 19107 16612 19156 16640
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 21082 16640 21088 16652
rect 19475 16612 21088 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21818 16600 21824 16652
rect 21876 16600 21882 16652
rect 21910 16600 21916 16652
rect 21968 16640 21974 16652
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 21968 16612 22385 16640
rect 21968 16600 21974 16612
rect 22373 16609 22385 16612
rect 22419 16609 22431 16643
rect 22373 16603 22431 16609
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 19242 16572 19248 16584
rect 18524 16544 19248 16572
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 21836 16572 21864 16600
rect 21836 16544 22094 16572
rect 16040 16476 16436 16504
rect 19705 16507 19763 16513
rect 19705 16473 19717 16507
rect 19751 16504 19763 16507
rect 19794 16504 19800 16516
rect 19751 16476 19800 16504
rect 19751 16473 19763 16476
rect 19705 16467 19763 16473
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 20438 16464 20444 16516
rect 20496 16464 20502 16516
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21453 16507 21511 16513
rect 21453 16504 21465 16507
rect 21324 16476 21465 16504
rect 21324 16464 21330 16476
rect 21453 16473 21465 16476
rect 21499 16473 21511 16507
rect 21453 16467 21511 16473
rect 5442 16436 5448 16448
rect 2746 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6454 16396 6460 16448
rect 6512 16436 6518 16448
rect 6641 16439 6699 16445
rect 6641 16436 6653 16439
rect 6512 16408 6653 16436
rect 6512 16396 6518 16408
rect 6641 16405 6653 16408
rect 6687 16405 6699 16439
rect 6641 16399 6699 16405
rect 7009 16439 7067 16445
rect 7009 16405 7021 16439
rect 7055 16436 7067 16439
rect 7558 16436 7564 16448
rect 7055 16408 7564 16436
rect 7055 16405 7067 16408
rect 7009 16399 7067 16405
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 7708 16408 7849 16436
rect 7708 16396 7714 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9214 16436 9220 16448
rect 9171 16408 9220 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11333 16439 11391 16445
rect 11333 16436 11345 16439
rect 11112 16408 11345 16436
rect 11112 16396 11118 16408
rect 11333 16405 11345 16408
rect 11379 16405 11391 16439
rect 11333 16399 11391 16405
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 13357 16439 13415 16445
rect 13357 16436 13369 16439
rect 12676 16408 13369 16436
rect 12676 16396 12682 16408
rect 13357 16405 13369 16408
rect 13403 16405 13415 16439
rect 13357 16399 13415 16405
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 15470 16396 15476 16448
rect 15528 16396 15534 16448
rect 17313 16439 17371 16445
rect 17313 16405 17325 16439
rect 17359 16436 17371 16439
rect 17402 16436 17408 16448
rect 17359 16408 17408 16436
rect 17359 16405 17371 16408
rect 17313 16399 17371 16405
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 18414 16396 18420 16448
rect 18472 16396 18478 16448
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 21913 16439 21971 16445
rect 21913 16436 21925 16439
rect 19116 16408 21925 16436
rect 19116 16396 19122 16408
rect 21913 16405 21925 16408
rect 21959 16405 21971 16439
rect 22066 16436 22094 16544
rect 22278 16532 22284 16584
rect 22336 16572 22342 16584
rect 22480 16572 22508 16603
rect 23934 16600 23940 16652
rect 23992 16600 23998 16652
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24946 16640 24952 16652
rect 24535 16612 24952 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 24946 16600 24952 16612
rect 25004 16640 25010 16652
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 25004 16612 25237 16640
rect 25004 16600 25010 16612
rect 25225 16609 25237 16612
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 25409 16643 25467 16649
rect 25409 16609 25421 16643
rect 25455 16640 25467 16643
rect 25682 16640 25688 16652
rect 25455 16612 25688 16640
rect 25455 16609 25467 16612
rect 25409 16603 25467 16609
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16640 26019 16643
rect 26050 16640 26056 16652
rect 26007 16612 26056 16640
rect 26007 16609 26019 16612
rect 25961 16603 26019 16609
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 26252 16649 26280 16680
rect 27724 16680 29736 16708
rect 27724 16649 27752 16680
rect 29730 16668 29736 16680
rect 29788 16668 29794 16720
rect 29840 16708 29868 16748
rect 31478 16708 31484 16720
rect 29840 16680 31484 16708
rect 26237 16643 26295 16649
rect 26237 16609 26249 16643
rect 26283 16609 26295 16643
rect 26237 16603 26295 16609
rect 27709 16643 27767 16649
rect 27709 16609 27721 16643
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 27798 16600 27804 16652
rect 27856 16600 27862 16652
rect 28718 16600 28724 16652
rect 28776 16640 28782 16652
rect 28905 16643 28963 16649
rect 28905 16640 28917 16643
rect 28776 16612 28917 16640
rect 28776 16600 28782 16612
rect 28905 16609 28917 16612
rect 28951 16609 28963 16643
rect 28905 16603 28963 16609
rect 29089 16643 29147 16649
rect 29089 16609 29101 16643
rect 29135 16640 29147 16643
rect 29840 16640 29868 16680
rect 31478 16668 31484 16680
rect 31536 16668 31542 16720
rect 29135 16612 29868 16640
rect 29135 16609 29147 16612
rect 29089 16603 29147 16609
rect 30006 16600 30012 16652
rect 30064 16600 30070 16652
rect 22336 16544 22508 16572
rect 23661 16575 23719 16581
rect 22336 16532 22342 16544
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 23750 16572 23756 16584
rect 23707 16544 23756 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16572 25191 16575
rect 26418 16572 26424 16584
rect 25179 16544 26424 16572
rect 25179 16541 25191 16544
rect 25133 16535 25191 16541
rect 23014 16464 23020 16516
rect 23072 16504 23078 16516
rect 25148 16504 25176 16535
rect 26418 16532 26424 16544
rect 26476 16532 26482 16584
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 28813 16575 28871 16581
rect 28813 16572 28825 16575
rect 27304 16544 28825 16572
rect 27304 16532 27310 16544
rect 28813 16541 28825 16544
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 29546 16532 29552 16584
rect 29604 16572 29610 16584
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29604 16544 29745 16572
rect 29604 16532 29610 16544
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 23072 16476 25176 16504
rect 23072 16464 23078 16476
rect 25314 16464 25320 16516
rect 25372 16504 25378 16516
rect 27617 16507 27675 16513
rect 25372 16476 27384 16504
rect 25372 16464 25378 16476
rect 22186 16436 22192 16448
rect 22066 16408 22192 16436
rect 21913 16399 21971 16405
rect 22186 16396 22192 16408
rect 22244 16436 22250 16448
rect 22281 16439 22339 16445
rect 22281 16436 22293 16439
rect 22244 16408 22293 16436
rect 22244 16396 22250 16408
rect 22281 16405 22293 16408
rect 22327 16405 22339 16439
rect 22281 16399 22339 16405
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 23198 16436 23204 16448
rect 22704 16408 23204 16436
rect 22704 16396 22710 16408
rect 23198 16396 23204 16408
rect 23256 16436 23262 16448
rect 23658 16436 23664 16448
rect 23256 16408 23664 16436
rect 23256 16396 23262 16408
rect 23658 16396 23664 16408
rect 23716 16436 23722 16448
rect 23753 16439 23811 16445
rect 23753 16436 23765 16439
rect 23716 16408 23765 16436
rect 23716 16396 23722 16408
rect 23753 16405 23765 16408
rect 23799 16405 23811 16439
rect 23753 16399 23811 16405
rect 24762 16396 24768 16448
rect 24820 16396 24826 16448
rect 27246 16396 27252 16448
rect 27304 16396 27310 16448
rect 27356 16436 27384 16476
rect 27617 16473 27629 16507
rect 27663 16504 27675 16507
rect 29362 16504 29368 16516
rect 27663 16476 29368 16504
rect 27663 16473 27675 16476
rect 27617 16467 27675 16473
rect 29362 16464 29368 16476
rect 29420 16464 29426 16516
rect 28445 16439 28503 16445
rect 28445 16436 28457 16439
rect 27356 16408 28457 16436
rect 28445 16405 28457 16408
rect 28491 16405 28503 16439
rect 28445 16399 28503 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 474 16192 480 16244
rect 532 16232 538 16244
rect 1118 16232 1124 16244
rect 532 16204 1124 16232
rect 532 16192 538 16204
rect 1118 16192 1124 16204
rect 1176 16192 1182 16244
rect 3786 16192 3792 16244
rect 3844 16232 3850 16244
rect 3844 16204 5580 16232
rect 3844 16192 3850 16204
rect 4430 16124 4436 16176
rect 4488 16124 4494 16176
rect 5552 16164 5580 16204
rect 5626 16192 5632 16244
rect 5684 16192 5690 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 6546 16232 6552 16244
rect 5767 16204 6552 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 8662 16232 8668 16244
rect 7883 16204 8668 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 8846 16192 8852 16244
rect 8904 16192 8910 16244
rect 8938 16192 8944 16244
rect 8996 16192 9002 16244
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 9456 16204 14841 16232
rect 9456 16192 9462 16204
rect 14829 16201 14841 16204
rect 14875 16201 14887 16235
rect 14829 16195 14887 16201
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 16540 16204 16681 16232
rect 16540 16192 16546 16204
rect 16669 16201 16681 16204
rect 16715 16201 16727 16235
rect 16669 16195 16727 16201
rect 16945 16235 17003 16241
rect 16945 16201 16957 16235
rect 16991 16232 17003 16235
rect 17034 16232 17040 16244
rect 16991 16204 17040 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 17034 16192 17040 16204
rect 17092 16232 17098 16244
rect 17865 16235 17923 16241
rect 17092 16204 17264 16232
rect 17092 16192 17098 16204
rect 7101 16167 7159 16173
rect 7101 16164 7113 16167
rect 5552 16136 7113 16164
rect 7101 16133 7113 16136
rect 7147 16133 7159 16167
rect 7101 16127 7159 16133
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 3326 16096 3332 16108
rect 1811 16068 3332 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3651 16068 6592 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 5905 16031 5963 16037
rect 5905 16028 5917 16031
rect 4856 16000 5917 16028
rect 4856 15988 4862 16000
rect 5905 15997 5917 16000
rect 5951 16028 5963 16031
rect 6362 16028 6368 16040
rect 5951 16000 6368 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 6564 15960 6592 16068
rect 7006 16056 7012 16108
rect 7064 16056 7070 16108
rect 7116 16096 7144 16127
rect 8386 16124 8392 16176
rect 8444 16164 8450 16176
rect 8864 16164 8892 16192
rect 9677 16167 9735 16173
rect 8444 16136 9260 16164
rect 8444 16124 8450 16136
rect 8570 16096 8576 16108
rect 7116 16068 8576 16096
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 9232 16096 9260 16136
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 9723 16136 10456 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 9140 16068 9260 16096
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 7650 16028 7656 16040
rect 7331 16000 7656 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 7742 15988 7748 16040
rect 7800 16028 7806 16040
rect 8662 16028 8668 16040
rect 7800 16000 8668 16028
rect 7800 15988 7806 16000
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 9140 16037 9168 16068
rect 9398 16056 9404 16108
rect 9456 16096 9462 16108
rect 9861 16099 9919 16105
rect 9456 16068 9674 16096
rect 9456 16056 9462 16068
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 15997 9183 16031
rect 9646 16028 9674 16068
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10134 16096 10140 16108
rect 9907 16068 10140 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10134 16056 10140 16068
rect 10192 16056 10198 16108
rect 10428 16096 10456 16136
rect 10502 16124 10508 16176
rect 10560 16124 10566 16176
rect 11333 16167 11391 16173
rect 11333 16133 11345 16167
rect 11379 16164 11391 16167
rect 12250 16164 12256 16176
rect 11379 16136 12256 16164
rect 11379 16133 11391 16136
rect 11333 16127 11391 16133
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 13814 16164 13820 16176
rect 13202 16136 13820 16164
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 14001 16167 14059 16173
rect 14001 16133 14013 16167
rect 14047 16164 14059 16167
rect 14090 16164 14096 16176
rect 14047 16136 14096 16164
rect 14047 16133 14059 16136
rect 14001 16127 14059 16133
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 17236 16164 17264 16204
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 19058 16232 19064 16244
rect 17911 16204 19064 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 19058 16192 19064 16204
rect 19116 16192 19122 16244
rect 20073 16235 20131 16241
rect 20073 16201 20085 16235
rect 20119 16232 20131 16235
rect 22465 16235 22523 16241
rect 20119 16204 22094 16232
rect 20119 16201 20131 16204
rect 20073 16195 20131 16201
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 14424 16136 17172 16164
rect 17236 16136 18521 16164
rect 14424 16124 14430 16136
rect 10870 16096 10876 16108
rect 10428 16068 10876 16096
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 14642 16096 14648 16108
rect 13320 16068 14648 16096
rect 13320 16056 13326 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15286 16096 15292 16108
rect 14967 16068 15292 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 9646 16000 10272 16028
rect 9125 15991 9183 15997
rect 7926 15960 7932 15972
rect 6564 15932 7932 15960
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 8478 15920 8484 15972
rect 8536 15920 8542 15972
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 9324 15932 10149 15960
rect 5261 15895 5319 15901
rect 5261 15861 5273 15895
rect 5307 15892 5319 15895
rect 6546 15892 6552 15904
rect 5307 15864 6552 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6638 15852 6644 15904
rect 6696 15852 6702 15904
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 9324 15892 9352 15932
rect 10137 15929 10149 15932
rect 10183 15929 10195 15963
rect 10244 15960 10272 16000
rect 10594 15988 10600 16040
rect 10652 15988 10658 16040
rect 10686 15988 10692 16040
rect 10744 15988 10750 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 10796 16000 11989 16028
rect 10796 15960 10824 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 14090 16028 14096 16040
rect 13044 16000 14096 16028
rect 13044 15988 13050 16000
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 15672 16028 15700 16059
rect 16022 16056 16028 16108
rect 16080 16096 16086 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16080 16068 17049 16096
rect 16080 16056 16086 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17144 16096 17172 16136
rect 18509 16133 18521 16136
rect 18555 16164 18567 16167
rect 18693 16167 18751 16173
rect 18693 16164 18705 16167
rect 18555 16136 18705 16164
rect 18555 16133 18567 16136
rect 18509 16127 18567 16133
rect 18693 16133 18705 16136
rect 18739 16164 18751 16167
rect 19426 16164 19432 16176
rect 18739 16136 19432 16164
rect 18739 16133 18751 16136
rect 18693 16127 18751 16133
rect 19426 16124 19432 16136
rect 19484 16164 19490 16176
rect 20530 16164 20536 16176
rect 19484 16136 20536 16164
rect 19484 16124 19490 16136
rect 20530 16124 20536 16136
rect 20588 16124 20594 16176
rect 22066 16164 22094 16204
rect 22465 16201 22477 16235
rect 22511 16232 22523 16235
rect 23290 16232 23296 16244
rect 22511 16204 23296 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 24121 16235 24179 16241
rect 24121 16201 24133 16235
rect 24167 16232 24179 16235
rect 27246 16232 27252 16244
rect 24167 16204 27252 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 24029 16167 24087 16173
rect 24029 16164 24041 16167
rect 22066 16136 24041 16164
rect 24029 16133 24041 16136
rect 24075 16133 24087 16167
rect 24029 16127 24087 16133
rect 26418 16124 26424 16176
rect 26476 16164 26482 16176
rect 27798 16164 27804 16176
rect 26476 16136 27804 16164
rect 26476 16124 26482 16136
rect 27798 16124 27804 16136
rect 27856 16164 27862 16176
rect 43530 16164 43536 16176
rect 27856 16136 43536 16164
rect 27856 16124 27862 16136
rect 43530 16124 43536 16136
rect 43588 16124 43594 16176
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 17144 16068 17785 16096
rect 17037 16059 17095 16065
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 19058 16096 19064 16108
rect 19015 16068 19064 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20438 16056 20444 16108
rect 20496 16056 20502 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 21542 16096 21548 16108
rect 21499 16068 21548 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 21542 16056 21548 16068
rect 21600 16056 21606 16108
rect 22557 16099 22615 16105
rect 22557 16065 22569 16099
rect 22603 16096 22615 16099
rect 23566 16096 23572 16108
rect 22603 16068 23572 16096
rect 22603 16065 22615 16068
rect 22557 16059 22615 16065
rect 23566 16056 23572 16068
rect 23624 16056 23630 16108
rect 26510 16096 26516 16108
rect 26266 16068 26516 16096
rect 26510 16056 26516 16068
rect 26568 16056 26574 16108
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27522 16096 27528 16108
rect 27212 16068 27528 16096
rect 27212 16056 27218 16068
rect 27522 16056 27528 16068
rect 27580 16056 27586 16108
rect 28261 16099 28319 16105
rect 28261 16065 28273 16099
rect 28307 16096 28319 16099
rect 28902 16096 28908 16108
rect 28307 16068 28908 16096
rect 28307 16065 28319 16068
rect 28261 16059 28319 16065
rect 28902 16056 28908 16068
rect 28960 16056 28966 16108
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 15672 16000 18061 16028
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 18598 16028 18604 16040
rect 18095 16000 18604 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 20530 15988 20536 16040
rect 20588 15988 20594 16040
rect 20625 16031 20683 16037
rect 20625 15997 20637 16031
rect 20671 16028 20683 16031
rect 22462 16028 22468 16040
rect 20671 16000 22468 16028
rect 20671 15997 20683 16000
rect 20625 15991 20683 15997
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 10244 15932 10824 15960
rect 10137 15923 10195 15929
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 15654 15960 15660 15972
rect 13688 15932 15660 15960
rect 13688 15920 13694 15932
rect 15654 15920 15660 15932
rect 15712 15960 15718 15972
rect 18506 15960 18512 15972
rect 15712 15932 18512 15960
rect 15712 15920 15718 15932
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 18782 15920 18788 15972
rect 18840 15960 18846 15972
rect 18966 15960 18972 15972
rect 18840 15932 18972 15960
rect 18840 15920 18846 15932
rect 18966 15920 18972 15932
rect 19024 15920 19030 15972
rect 20162 15920 20168 15972
rect 20220 15960 20226 15972
rect 22097 15963 22155 15969
rect 22097 15960 22109 15963
rect 20220 15932 22109 15960
rect 20220 15920 20226 15932
rect 22097 15929 22109 15932
rect 22143 15929 22155 15963
rect 22097 15923 22155 15929
rect 8628 15864 9352 15892
rect 8628 15852 8634 15864
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 9858 15892 9864 15904
rect 9548 15864 9864 15892
rect 9548 15852 9554 15864
rect 9858 15852 9864 15864
rect 9916 15892 9922 15904
rect 10594 15892 10600 15904
rect 9916 15864 10600 15892
rect 9916 15852 9922 15864
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11606 15892 11612 15904
rect 11112 15864 11612 15892
rect 11112 15852 11118 15864
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 11974 15892 11980 15904
rect 11848 15864 11980 15892
rect 11848 15852 11854 15864
rect 11974 15852 11980 15864
rect 12032 15892 12038 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12032 15864 13461 15892
rect 12032 15852 12038 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 13814 15852 13820 15904
rect 13872 15852 13878 15904
rect 14461 15895 14519 15901
rect 14461 15861 14473 15895
rect 14507 15892 14519 15895
rect 16022 15892 16028 15904
rect 14507 15864 16028 15892
rect 14507 15861 14519 15864
rect 14461 15855 14519 15861
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16482 15892 16488 15904
rect 16347 15864 16488 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 17368 15864 17417 15892
rect 17368 15852 17374 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 19610 15852 19616 15904
rect 19668 15852 19674 15904
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 20772 15864 21281 15892
rect 20772 15852 20778 15864
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21269 15855 21327 15861
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 22664 15892 22692 15991
rect 23198 15988 23204 16040
rect 23256 16028 23262 16040
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 23256 16000 23305 16028
rect 23256 15988 23262 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 24305 16031 24363 16037
rect 24305 15997 24317 16031
rect 24351 15997 24363 16031
rect 24305 15991 24363 15997
rect 22738 15920 22744 15972
rect 22796 15960 22802 15972
rect 23661 15963 23719 15969
rect 23661 15960 23673 15963
rect 22796 15932 23673 15960
rect 22796 15920 22802 15932
rect 23661 15929 23673 15932
rect 23707 15929 23719 15963
rect 23661 15923 23719 15929
rect 21784 15864 22692 15892
rect 23201 15895 23259 15901
rect 21784 15852 21790 15864
rect 23201 15861 23213 15895
rect 23247 15892 23259 15895
rect 23566 15892 23572 15904
rect 23247 15864 23572 15892
rect 23247 15861 23259 15864
rect 23201 15855 23259 15861
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 24320 15892 24348 15991
rect 24854 15988 24860 16040
rect 24912 15988 24918 16040
rect 25133 16031 25191 16037
rect 25133 15997 25145 16031
rect 25179 16028 25191 16031
rect 27801 16031 27859 16037
rect 27801 16028 27813 16031
rect 25179 16000 27813 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27801 15997 27813 16000
rect 27847 15997 27859 16031
rect 27801 15991 27859 15997
rect 26142 15920 26148 15972
rect 26200 15960 26206 15972
rect 28905 15963 28963 15969
rect 28905 15960 28917 15963
rect 26200 15932 28917 15960
rect 26200 15920 26206 15932
rect 28905 15929 28917 15932
rect 28951 15929 28963 15963
rect 28905 15923 28963 15929
rect 29012 15932 29684 15960
rect 26605 15895 26663 15901
rect 26605 15892 26617 15895
rect 24320 15864 26617 15892
rect 26605 15861 26617 15864
rect 26651 15892 26663 15895
rect 27614 15892 27620 15904
rect 26651 15864 27620 15892
rect 26651 15861 26663 15864
rect 26605 15855 26663 15861
rect 27614 15852 27620 15864
rect 27672 15852 27678 15904
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 29012 15892 29040 15932
rect 27764 15864 29040 15892
rect 27764 15852 27770 15864
rect 29546 15852 29552 15904
rect 29604 15852 29610 15904
rect 29656 15892 29684 15932
rect 30374 15920 30380 15972
rect 30432 15960 30438 15972
rect 46934 15960 46940 15972
rect 30432 15932 46940 15960
rect 30432 15920 30438 15932
rect 46934 15920 46940 15932
rect 46992 15920 46998 15972
rect 45278 15892 45284 15904
rect 29656 15864 45284 15892
rect 45278 15852 45284 15864
rect 45336 15852 45342 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 5684 15660 6868 15688
rect 5684 15648 5690 15660
rect 5169 15623 5227 15629
rect 5169 15589 5181 15623
rect 5215 15620 5227 15623
rect 6730 15620 6736 15632
rect 5215 15592 6736 15620
rect 5215 15589 5227 15592
rect 5169 15583 5227 15589
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 6840 15620 6868 15660
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7616 15660 7849 15688
rect 7616 15648 7622 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 9398 15688 9404 15700
rect 7984 15660 9404 15688
rect 7984 15648 7990 15660
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9628 15648 9634 15700
rect 9686 15688 9692 15700
rect 10502 15688 10508 15700
rect 9686 15660 10508 15688
rect 9686 15648 9692 15660
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 13265 15691 13323 15697
rect 10652 15660 12112 15688
rect 10652 15648 10658 15660
rect 7469 15623 7527 15629
rect 6840 15592 6960 15620
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4890 15552 4896 15564
rect 4663 15524 4896 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 6362 15552 6368 15564
rect 5859 15524 6368 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 6932 15561 6960 15592
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 8754 15620 8760 15632
rect 7515 15592 8760 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9766 15620 9772 15632
rect 8864 15592 9772 15620
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6604 15524 6837 15552
rect 6604 15512 6610 15524
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 8478 15512 8484 15564
rect 8536 15512 8542 15564
rect 8662 15512 8668 15564
rect 8720 15552 8726 15564
rect 8864 15552 8892 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 11422 15580 11428 15632
rect 11480 15620 11486 15632
rect 12084 15620 12112 15660
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 13446 15688 13452 15700
rect 13311 15660 13452 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 15470 15688 15476 15700
rect 14783 15660 15476 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18877 15691 18935 15697
rect 18877 15688 18889 15691
rect 17828 15660 18889 15688
rect 17828 15648 17834 15660
rect 18877 15657 18889 15660
rect 18923 15657 18935 15691
rect 18877 15651 18935 15657
rect 18966 15648 18972 15700
rect 19024 15688 19030 15700
rect 19024 15660 24624 15688
rect 19024 15648 19030 15660
rect 20530 15620 20536 15632
rect 11480 15592 12020 15620
rect 12084 15592 17264 15620
rect 11480 15580 11486 15592
rect 8720 15524 8892 15552
rect 8720 15512 8726 15524
rect 9628 15512 9634 15564
rect 9686 15552 9692 15564
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 9686 15524 10149 15552
rect 9686 15512 9692 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10318 15512 10324 15564
rect 10376 15512 10382 15564
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 10652 15524 11529 15552
rect 10652 15512 10658 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 11992 15552 12020 15592
rect 12805 15555 12863 15561
rect 11992 15524 12756 15552
rect 11517 15515 11575 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 3510 15484 3516 15496
rect 1811 15456 3516 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 4246 15444 4252 15496
rect 4304 15484 4310 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4304 15456 4445 15484
rect 4304 15444 4310 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 5534 15444 5540 15496
rect 5592 15444 5598 15496
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 7834 15484 7840 15496
rect 6779 15456 7840 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 7926 15444 7932 15496
rect 7984 15484 7990 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 7984 15456 9229 15484
rect 7984 15444 7990 15456
rect 9217 15453 9229 15456
rect 9263 15484 9275 15487
rect 9858 15484 9864 15496
rect 9263 15456 9864 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10410 15484 10416 15496
rect 10091 15456 10416 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15484 11391 15487
rect 11606 15484 11612 15496
rect 11379 15456 11612 15484
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 11992 15456 12541 15484
rect 5629 15419 5687 15425
rect 5629 15416 5641 15419
rect 3988 15388 5641 15416
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 2740 15320 3341 15348
rect 2740 15308 2746 15320
rect 3329 15317 3341 15320
rect 3375 15348 3387 15351
rect 3513 15351 3571 15357
rect 3513 15348 3525 15351
rect 3375 15320 3525 15348
rect 3375 15317 3387 15320
rect 3329 15311 3387 15317
rect 3513 15317 3525 15320
rect 3559 15348 3571 15351
rect 3786 15348 3792 15360
rect 3559 15320 3792 15348
rect 3559 15317 3571 15320
rect 3513 15311 3571 15317
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 3988 15357 4016 15388
rect 5629 15385 5641 15388
rect 5675 15385 5687 15419
rect 5629 15379 5687 15385
rect 6454 15376 6460 15428
rect 6512 15416 6518 15428
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 6512 15388 8309 15416
rect 6512 15376 6518 15388
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 8662 15376 8668 15428
rect 8720 15416 8726 15428
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 8720 15388 9321 15416
rect 8720 15376 8726 15388
rect 9309 15385 9321 15388
rect 9355 15416 9367 15419
rect 9398 15416 9404 15428
rect 9355 15388 9404 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 9398 15376 9404 15388
rect 9456 15376 9462 15428
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 11422 15416 11428 15428
rect 9640 15388 11428 15416
rect 9640 15376 9646 15388
rect 11422 15376 11428 15388
rect 11480 15376 11486 15428
rect 3973 15351 4031 15357
rect 3973 15317 3985 15351
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 4338 15308 4344 15360
rect 4396 15308 4402 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 6365 15351 6423 15357
rect 6365 15348 6377 15351
rect 5500 15320 6377 15348
rect 5500 15308 5506 15320
rect 6365 15317 6377 15320
rect 6411 15317 6423 15351
rect 6365 15311 6423 15317
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7524 15320 8217 15348
rect 7524 15308 7530 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8205 15311 8263 15317
rect 8754 15308 8760 15360
rect 8812 15348 8818 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8812 15320 8953 15348
rect 8812 15308 8818 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 9916 15320 10977 15348
rect 9916 15308 9922 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11992 15357 12020 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12728 15484 12756 15524
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 13630 15552 13636 15564
rect 12851 15524 13636 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15552 14519 15555
rect 14826 15552 14832 15564
rect 14507 15524 14832 15552
rect 14507 15521 14519 15524
rect 14461 15515 14519 15521
rect 14826 15512 14832 15524
rect 14884 15552 14890 15564
rect 15197 15555 15255 15561
rect 15197 15552 15209 15555
rect 14884 15524 15209 15552
rect 14884 15512 14890 15524
rect 15197 15521 15209 15524
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 15654 15552 15660 15564
rect 15427 15524 15660 15552
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 15654 15512 15660 15524
rect 15712 15512 15718 15564
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16758 15552 16764 15564
rect 16623 15524 16764 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 16758 15512 16764 15524
rect 16816 15552 16822 15564
rect 16816 15524 17080 15552
rect 16816 15512 16822 15524
rect 13262 15484 13268 15496
rect 12728 15456 13268 15484
rect 12529 15447 12587 15453
rect 13262 15444 13268 15456
rect 13320 15444 13326 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 15562 15484 15568 15496
rect 13771 15456 15568 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16850 15484 16856 15496
rect 16439 15456 16856 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 14200 15388 15117 15416
rect 14200 15360 14228 15388
rect 15105 15385 15117 15388
rect 15151 15385 15163 15419
rect 15105 15379 15163 15385
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 16758 15416 16764 15428
rect 15252 15388 16764 15416
rect 15252 15376 15258 15388
rect 16758 15376 16764 15388
rect 16816 15376 16822 15428
rect 11977 15351 12035 15357
rect 11977 15348 11989 15351
rect 11572 15320 11989 15348
rect 11572 15308 11578 15320
rect 11977 15317 11989 15320
rect 12023 15317 12035 15351
rect 11977 15311 12035 15317
rect 12158 15308 12164 15360
rect 12216 15308 12222 15360
rect 12618 15308 12624 15360
rect 12676 15308 12682 15360
rect 13538 15308 13544 15360
rect 13596 15308 13602 15360
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 16206 15308 16212 15360
rect 16264 15348 16270 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16264 15320 16313 15348
rect 16264 15308 16270 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 17052 15348 17080 15524
rect 17126 15512 17132 15564
rect 17184 15512 17190 15564
rect 17236 15552 17264 15592
rect 18432 15592 20536 15620
rect 18432 15552 18460 15592
rect 20530 15580 20536 15592
rect 20588 15620 20594 15632
rect 20717 15623 20775 15629
rect 20717 15620 20729 15623
rect 20588 15592 20729 15620
rect 20588 15580 20594 15592
rect 20717 15589 20729 15592
rect 20763 15589 20775 15623
rect 20717 15583 20775 15589
rect 22462 15580 22468 15632
rect 22520 15620 22526 15632
rect 22520 15592 24532 15620
rect 22520 15580 22526 15592
rect 19337 15555 19395 15561
rect 19337 15552 19349 15555
rect 17236 15524 18460 15552
rect 18524 15524 19349 15552
rect 18524 15470 18552 15524
rect 19337 15521 19349 15524
rect 19383 15552 19395 15555
rect 19426 15552 19432 15564
rect 19383 15524 19432 15552
rect 19383 15521 19395 15524
rect 19337 15515 19395 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 20162 15512 20168 15564
rect 20220 15512 20226 15564
rect 20349 15555 20407 15561
rect 20349 15521 20361 15555
rect 20395 15552 20407 15555
rect 20990 15552 20996 15564
rect 20395 15524 20996 15552
rect 20395 15521 20407 15524
rect 20349 15515 20407 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 22094 15552 22100 15564
rect 21140 15524 22100 15552
rect 21140 15512 21146 15524
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 23842 15512 23848 15564
rect 23900 15512 23906 15564
rect 24504 15484 24532 15592
rect 24596 15561 24624 15660
rect 26602 15648 26608 15700
rect 26660 15688 26666 15700
rect 26660 15660 27016 15688
rect 26660 15648 26666 15660
rect 24946 15580 24952 15632
rect 25004 15620 25010 15632
rect 25004 15592 26924 15620
rect 25004 15580 25010 15592
rect 26896 15564 26924 15592
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 25740 15524 25789 15552
rect 25740 15512 25746 15524
rect 25777 15521 25789 15524
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 26878 15512 26884 15564
rect 26936 15512 26942 15564
rect 26988 15561 27016 15660
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 28629 15691 28687 15697
rect 28629 15688 28641 15691
rect 28592 15660 28641 15688
rect 28592 15648 28598 15660
rect 28629 15657 28641 15660
rect 28675 15688 28687 15691
rect 28718 15688 28724 15700
rect 28675 15660 28724 15688
rect 28675 15657 28687 15660
rect 28629 15651 28687 15657
rect 28718 15648 28724 15660
rect 28776 15648 28782 15700
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 27154 15484 27160 15496
rect 24504 15456 27160 15484
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27614 15444 27620 15496
rect 27672 15444 27678 15496
rect 17402 15376 17408 15428
rect 17460 15376 17466 15428
rect 18966 15376 18972 15428
rect 19024 15416 19030 15428
rect 19024 15388 20208 15416
rect 19024 15376 19030 15388
rect 18874 15348 18880 15360
rect 17052 15320 18880 15348
rect 16301 15311 16359 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19242 15308 19248 15360
rect 19300 15348 19306 15360
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 19300 15320 19717 15348
rect 19300 15308 19306 15320
rect 19705 15317 19717 15320
rect 19751 15317 19763 15351
rect 19705 15311 19763 15317
rect 20070 15308 20076 15360
rect 20128 15308 20134 15360
rect 20180 15348 20208 15388
rect 20622 15376 20628 15428
rect 20680 15416 20686 15428
rect 21082 15416 21088 15428
rect 20680 15388 21088 15416
rect 20680 15376 20686 15388
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 21358 15376 21364 15428
rect 21416 15376 21422 15428
rect 23566 15416 23572 15428
rect 22586 15388 23572 15416
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 23658 15376 23664 15428
rect 23716 15416 23722 15428
rect 24302 15416 24308 15428
rect 23716 15388 24308 15416
rect 23716 15376 23722 15388
rect 24302 15376 24308 15388
rect 24360 15376 24366 15428
rect 25685 15419 25743 15425
rect 25685 15385 25697 15419
rect 25731 15416 25743 15419
rect 26142 15416 26148 15428
rect 25731 15388 26148 15416
rect 25731 15385 25743 15388
rect 25685 15379 25743 15385
rect 26142 15376 26148 15388
rect 26200 15376 26206 15428
rect 26789 15419 26847 15425
rect 26789 15385 26801 15419
rect 26835 15416 26847 15419
rect 27798 15416 27804 15428
rect 26835 15388 27804 15416
rect 26835 15385 26847 15388
rect 26789 15379 26847 15385
rect 27798 15376 27804 15388
rect 27856 15376 27862 15428
rect 21726 15348 21732 15360
rect 20180 15320 21732 15348
rect 21726 15308 21732 15320
rect 21784 15348 21790 15360
rect 22833 15351 22891 15357
rect 22833 15348 22845 15351
rect 21784 15320 22845 15348
rect 21784 15308 21790 15320
rect 22833 15317 22845 15320
rect 22879 15317 22891 15351
rect 22833 15311 22891 15317
rect 23290 15308 23296 15360
rect 23348 15308 23354 15360
rect 23753 15351 23811 15357
rect 23753 15317 23765 15351
rect 23799 15348 23811 15351
rect 24394 15348 24400 15360
rect 23799 15320 24400 15348
rect 23799 15317 23811 15320
rect 23753 15311 23811 15317
rect 24394 15308 24400 15320
rect 24452 15308 24458 15360
rect 25222 15308 25228 15360
rect 25280 15308 25286 15360
rect 25590 15308 25596 15360
rect 25648 15308 25654 15360
rect 25774 15308 25780 15360
rect 25832 15348 25838 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 25832 15320 26433 15348
rect 25832 15308 25838 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 26421 15311 26479 15317
rect 26970 15308 26976 15360
rect 27028 15348 27034 15360
rect 28261 15351 28319 15357
rect 28261 15348 28273 15351
rect 27028 15320 28273 15348
rect 27028 15308 27034 15320
rect 28261 15317 28273 15320
rect 28307 15317 28319 15351
rect 28261 15311 28319 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 198 15104 204 15156
rect 256 15144 262 15156
rect 1118 15144 1124 15156
rect 256 15116 1124 15144
rect 256 15104 262 15116
rect 1118 15104 1124 15116
rect 1176 15104 1182 15156
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 4982 15104 4988 15156
rect 5040 15104 5046 15156
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 7834 15144 7840 15156
rect 6604 15116 7840 15144
rect 6604 15104 6610 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8478 15144 8484 15156
rect 8260 15116 8484 15144
rect 8260 15104 8266 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8588 15116 12388 15144
rect 8588 15076 8616 15116
rect 3528 15048 8616 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 3418 15008 3424 15020
rect 1811 14980 3424 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 3528 15017 3556 15048
rect 8754 15036 8760 15088
rect 8812 15036 8818 15088
rect 9490 15036 9496 15088
rect 9548 15076 9554 15088
rect 9548 15048 9812 15076
rect 9548 15036 9554 15048
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6362 15008 6368 15020
rect 6236 14980 6368 15008
rect 6236 14968 6242 14980
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 1118 14900 1124 14952
rect 1176 14940 1182 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1176 14912 2053 14940
rect 1176 14900 1182 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 4212 14912 5089 14940
rect 4212 14900 4218 14912
rect 5077 14909 5089 14912
rect 5123 14909 5135 14943
rect 5077 14903 5135 14909
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5626 14940 5632 14952
rect 5307 14912 5632 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 6840 14940 6868 14971
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 6972 14980 7941 15008
rect 6972 14968 6978 14980
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 9784 15008 9812 15048
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10134 15076 10140 15088
rect 10008 15048 10140 15076
rect 10008 15036 10014 15048
rect 10134 15036 10140 15048
rect 10192 15036 10198 15088
rect 12360 15076 12388 15116
rect 12434 15104 12440 15156
rect 12492 15104 12498 15156
rect 16298 15104 16304 15156
rect 16356 15104 16362 15156
rect 17034 15104 17040 15156
rect 17092 15104 17098 15156
rect 18230 15104 18236 15156
rect 18288 15144 18294 15156
rect 19518 15144 19524 15156
rect 18288 15116 19524 15144
rect 18288 15104 18294 15116
rect 19518 15104 19524 15116
rect 19576 15144 19582 15156
rect 20622 15144 20628 15156
rect 19576 15116 20628 15144
rect 19576 15104 19582 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 21266 15144 21272 15156
rect 20772 15116 21272 15144
rect 20772 15104 20778 15116
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 21358 15104 21364 15156
rect 21416 15144 21422 15156
rect 27154 15144 27160 15156
rect 21416 15116 27160 15144
rect 21416 15104 21422 15116
rect 27154 15104 27160 15116
rect 27212 15104 27218 15156
rect 27430 15104 27436 15156
rect 27488 15104 27494 15156
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 27798 15144 27804 15156
rect 27663 15116 27804 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 27798 15104 27804 15116
rect 27856 15104 27862 15156
rect 10244 15048 11008 15076
rect 12360 15048 12756 15076
rect 10244 15008 10272 15048
rect 9784 14980 10272 15008
rect 7929 14971 7987 14977
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10744 14980 10793 15008
rect 10744 14968 10750 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 7742 14940 7748 14952
rect 6840 14912 7748 14940
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 10594 14940 10600 14952
rect 8260 14912 9352 14940
rect 8260 14900 8266 14912
rect 6549 14875 6607 14881
rect 6549 14841 6561 14875
rect 6595 14872 6607 14875
rect 9324 14872 9352 14912
rect 9508 14912 10600 14940
rect 9508 14872 9536 14912
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10980 14949 11008 15048
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11664 14980 11805 15008
rect 11664 14968 11670 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14909 11023 14943
rect 12728 14940 12756 15048
rect 13262 15036 13268 15088
rect 13320 15076 13326 15088
rect 14829 15079 14887 15085
rect 14829 15076 14841 15079
rect 13320 15048 14841 15076
rect 13320 15036 13326 15048
rect 14829 15045 14841 15048
rect 14875 15045 14887 15079
rect 14829 15039 14887 15045
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 19334 15076 19340 15088
rect 16448 15048 19340 15076
rect 16448 15036 16454 15048
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 19610 15036 19616 15088
rect 19668 15076 19674 15088
rect 19981 15079 20039 15085
rect 19981 15076 19993 15079
rect 19668 15048 19993 15076
rect 19668 15036 19674 15048
rect 19981 15045 19993 15048
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 20530 15036 20536 15088
rect 20588 15036 20594 15088
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 23845 15079 23903 15085
rect 23845 15076 23857 15079
rect 22152 15048 23857 15076
rect 22152 15036 22158 15048
rect 23845 15045 23857 15048
rect 23891 15076 23903 15079
rect 24854 15076 24860 15088
rect 23891 15048 24860 15076
rect 23891 15045 23903 15048
rect 23845 15039 23903 15045
rect 24854 15036 24860 15048
rect 24912 15036 24918 15088
rect 26878 15036 26884 15088
rect 26936 15076 26942 15088
rect 27709 15079 27767 15085
rect 27709 15076 27721 15079
rect 26936 15048 27721 15076
rect 26936 15036 26942 15048
rect 27709 15045 27721 15048
rect 27755 15076 27767 15079
rect 27755 15048 31754 15076
rect 27755 15045 27767 15048
rect 27709 15039 27767 15045
rect 12802 14968 12808 15020
rect 12860 14968 12866 15020
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 15008 12955 15011
rect 13538 15008 13544 15020
rect 12943 14980 13544 15008
rect 12943 14977 12955 14980
rect 12897 14971 12955 14977
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 16298 15008 16304 15020
rect 15962 14980 16304 15008
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 15008 17371 15011
rect 19426 15008 19432 15020
rect 17359 14980 19432 15008
rect 17359 14977 17371 14980
rect 17313 14971 17371 14977
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 19702 14968 19708 15020
rect 19760 14968 19766 15020
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 12989 14943 13047 14949
rect 12989 14940 13001 14943
rect 12728 14912 13001 14940
rect 10965 14903 11023 14909
rect 12989 14909 13001 14912
rect 13035 14940 13047 14943
rect 13722 14940 13728 14952
rect 13035 14912 13728 14940
rect 13035 14909 13047 14912
rect 12989 14903 13047 14909
rect 10888 14872 10916 14903
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 16206 14940 16212 14952
rect 13832 14912 16212 14940
rect 13832 14872 13860 14912
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16942 14940 16948 14952
rect 16316 14912 16948 14940
rect 6595 14844 8064 14872
rect 9324 14844 9536 14872
rect 9646 14844 12020 14872
rect 6595 14841 6607 14844
rect 6549 14835 6607 14841
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 5810 14764 5816 14816
rect 5868 14764 5874 14816
rect 7466 14764 7472 14816
rect 7524 14764 7530 14816
rect 8036 14804 8064 14844
rect 9646 14816 9674 14844
rect 8938 14804 8944 14816
rect 8036 14776 8944 14804
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9582 14764 9588 14816
rect 9640 14776 9674 14816
rect 9640 14764 9646 14776
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 10413 14807 10471 14813
rect 10413 14804 10425 14807
rect 10008 14776 10425 14804
rect 10008 14764 10014 14776
rect 10413 14773 10425 14776
rect 10459 14773 10471 14807
rect 10413 14767 10471 14773
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 10560 14776 11897 14804
rect 10560 14764 10566 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 11992 14804 12020 14844
rect 13372 14844 13860 14872
rect 13372 14804 13400 14844
rect 13906 14832 13912 14884
rect 13964 14832 13970 14884
rect 11992 14776 13400 14804
rect 11885 14767 11943 14773
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 16316 14804 16344 14912
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17402 14900 17408 14952
rect 17460 14940 17466 14952
rect 20714 14940 20720 14952
rect 17460 14912 20720 14940
rect 17460 14900 17466 14912
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 21453 14943 21511 14949
rect 21453 14940 21465 14943
rect 21048 14912 21465 14940
rect 21048 14900 21054 14912
rect 21453 14909 21465 14912
rect 21499 14940 21511 14943
rect 22020 14940 22048 14971
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 22520 14980 23121 15008
rect 22520 14968 22526 14980
rect 23109 14977 23121 14980
rect 23155 15008 23167 15011
rect 23382 15008 23388 15020
rect 23155 14980 23388 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 26510 15008 26516 15020
rect 26266 14980 26516 15008
rect 26510 14968 26516 14980
rect 26568 15008 26574 15020
rect 27430 15008 27436 15020
rect 26568 14980 27436 15008
rect 26568 14968 26574 14980
rect 27430 14968 27436 14980
rect 27488 14968 27494 15020
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 27893 15011 27951 15017
rect 27893 15008 27905 15011
rect 27672 14980 27905 15008
rect 27672 14968 27678 14980
rect 27893 14977 27905 14980
rect 27939 15008 27951 15011
rect 27939 14980 28994 15008
rect 27939 14977 27951 14980
rect 27893 14971 27951 14977
rect 21499 14912 22048 14940
rect 24857 14943 24915 14949
rect 21499 14909 21511 14912
rect 21453 14903 21511 14909
rect 24857 14909 24869 14943
rect 24903 14940 24915 14943
rect 25133 14943 25191 14949
rect 24903 14912 24992 14940
rect 24903 14909 24915 14912
rect 24857 14903 24915 14909
rect 16758 14832 16764 14884
rect 16816 14872 16822 14884
rect 18230 14872 18236 14884
rect 16816 14844 18236 14872
rect 16816 14832 16822 14844
rect 18230 14832 18236 14844
rect 18288 14872 18294 14884
rect 18601 14875 18659 14881
rect 18601 14872 18613 14875
rect 18288 14844 18613 14872
rect 18288 14832 18294 14844
rect 18601 14841 18613 14844
rect 18647 14841 18659 14875
rect 18601 14835 18659 14841
rect 18782 14832 18788 14884
rect 18840 14872 18846 14884
rect 19150 14872 19156 14884
rect 18840 14844 19156 14872
rect 18840 14832 18846 14844
rect 19150 14832 19156 14844
rect 19208 14872 19214 14884
rect 19208 14844 19840 14872
rect 19208 14832 19214 14844
rect 13596 14776 16344 14804
rect 13596 14764 13602 14776
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 19334 14804 19340 14816
rect 17000 14776 19340 14804
rect 17000 14764 17006 14776
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19426 14764 19432 14816
rect 19484 14764 19490 14816
rect 19812 14804 19840 14844
rect 21358 14832 21364 14884
rect 21416 14872 21422 14884
rect 21416 14844 24440 14872
rect 21416 14832 21422 14844
rect 24412 14816 24440 14844
rect 20990 14804 20996 14816
rect 19812 14776 20996 14804
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 22649 14807 22707 14813
rect 22649 14804 22661 14807
rect 22612 14776 22661 14804
rect 22612 14764 22618 14776
rect 22649 14773 22661 14776
rect 22695 14773 22707 14807
rect 22649 14767 22707 14773
rect 24302 14764 24308 14816
rect 24360 14764 24366 14816
rect 24394 14764 24400 14816
rect 24452 14804 24458 14816
rect 24581 14807 24639 14813
rect 24581 14804 24593 14807
rect 24452 14776 24593 14804
rect 24452 14764 24458 14776
rect 24581 14773 24593 14776
rect 24627 14804 24639 14807
rect 24854 14804 24860 14816
rect 24627 14776 24860 14804
rect 24627 14773 24639 14776
rect 24581 14767 24639 14773
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 24964 14804 24992 14912
rect 25133 14909 25145 14943
rect 25179 14940 25191 14943
rect 26970 14940 26976 14952
rect 25179 14912 26976 14940
rect 25179 14909 25191 14912
rect 25133 14903 25191 14909
rect 26970 14900 26976 14912
rect 27028 14900 27034 14952
rect 26142 14832 26148 14884
rect 26200 14872 26206 14884
rect 27249 14875 27307 14881
rect 27249 14872 27261 14875
rect 26200 14844 27261 14872
rect 26200 14832 26206 14844
rect 27249 14841 27261 14844
rect 27295 14872 27307 14875
rect 28966 14872 28994 14980
rect 31726 14940 31754 15048
rect 43438 14940 43444 14952
rect 31726 14912 43444 14940
rect 43438 14900 43444 14912
rect 43496 14900 43502 14952
rect 46198 14872 46204 14884
rect 27295 14844 28028 14872
rect 28966 14844 46204 14872
rect 27295 14841 27307 14844
rect 27249 14835 27307 14841
rect 25866 14804 25872 14816
rect 24964 14776 25872 14804
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 26234 14764 26240 14816
rect 26292 14804 26298 14816
rect 26602 14804 26608 14816
rect 26292 14776 26608 14804
rect 26292 14764 26298 14776
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 27065 14807 27123 14813
rect 27065 14773 27077 14807
rect 27111 14804 27123 14807
rect 27430 14804 27436 14816
rect 27111 14776 27436 14804
rect 27111 14773 27123 14776
rect 27065 14767 27123 14773
rect 27430 14764 27436 14776
rect 27488 14764 27494 14816
rect 28000 14804 28028 14844
rect 46198 14832 46204 14844
rect 46256 14832 46262 14884
rect 48590 14804 48596 14816
rect 28000 14776 48596 14804
rect 48590 14764 48596 14776
rect 48648 14764 48654 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 4154 14560 4160 14612
rect 4212 14560 4218 14612
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 8536 14572 9413 14600
rect 8536 14560 8542 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 9646 14572 9904 14600
rect 7650 14532 7656 14544
rect 6656 14504 7656 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 3602 14424 3608 14476
rect 3660 14424 3666 14476
rect 4798 14424 4804 14476
rect 4856 14424 4862 14476
rect 4890 14424 4896 14476
rect 4948 14464 4954 14476
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 4948 14436 5641 14464
rect 4948 14424 4954 14436
rect 5629 14433 5641 14436
rect 5675 14464 5687 14467
rect 6656 14464 6684 14504
rect 7650 14492 7656 14504
rect 7708 14532 7714 14544
rect 9214 14532 9220 14544
rect 7708 14504 9220 14532
rect 7708 14492 7714 14504
rect 5675 14436 6684 14464
rect 7377 14467 7435 14473
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 7558 14464 7564 14476
rect 7423 14436 7564 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 8404 14473 8432 14504
rect 9214 14492 9220 14504
rect 9272 14492 9278 14544
rect 9646 14532 9674 14572
rect 9324 14504 9674 14532
rect 8297 14467 8355 14473
rect 8297 14464 8309 14467
rect 8260 14436 8309 14464
rect 8260 14424 8266 14436
rect 8297 14433 8309 14436
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 5166 14396 5172 14408
rect 1811 14368 5172 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5350 14356 5356 14408
rect 5408 14356 5414 14408
rect 8312 14396 8340 14427
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 9324 14464 9352 14504
rect 9766 14492 9772 14544
rect 9824 14492 9830 14544
rect 9876 14532 9904 14572
rect 11698 14560 11704 14612
rect 11756 14560 11762 14612
rect 13722 14560 13728 14612
rect 13780 14560 13786 14612
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 14148 14572 14197 14600
rect 14148 14560 14154 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 17310 14600 17316 14612
rect 14185 14563 14243 14569
rect 14292 14572 17316 14600
rect 11974 14532 11980 14544
rect 9876 14504 11980 14532
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 14292 14532 14320 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 18564 14572 18613 14600
rect 18564 14560 18570 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 18690 14560 18696 14612
rect 18748 14600 18754 14612
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18748 14572 18981 14600
rect 18748 14560 18754 14572
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 13596 14504 14320 14532
rect 13596 14492 13602 14504
rect 9784 14464 9812 14492
rect 8536 14436 9352 14464
rect 9646 14436 9812 14464
rect 8536 14424 8542 14436
rect 9646 14396 9674 14436
rect 9858 14424 9864 14476
rect 9916 14424 9922 14476
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10134 14464 10140 14476
rect 10091 14436 10140 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10284 14436 11161 14464
rect 10284 14424 10290 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 14182 14464 14188 14476
rect 11149 14427 11207 14433
rect 11256 14436 14188 14464
rect 8312 14368 9674 14396
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 10594 14396 10600 14408
rect 9815 14368 10600 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 10928 14368 11069 14396
rect 10928 14356 10934 14368
rect 11057 14365 11069 14368
rect 11103 14396 11115 14399
rect 11256 14396 11284 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15378 14464 15384 14476
rect 14967 14436 15384 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 18414 14464 18420 14476
rect 17175 14436 18420 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 11103 14368 11284 14396
rect 11103 14365 11115 14368
rect 11057 14359 11115 14365
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 18984 14396 19012 14563
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 19978 14600 19984 14612
rect 19300 14572 19984 14600
rect 19300 14560 19306 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20622 14560 20628 14612
rect 20680 14600 20686 14612
rect 21818 14600 21824 14612
rect 20680 14572 21824 14600
rect 20680 14560 20686 14572
rect 21818 14560 21824 14572
rect 21876 14600 21882 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21876 14572 21925 14600
rect 21876 14560 21882 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 21913 14563 21971 14569
rect 24029 14603 24087 14609
rect 24029 14569 24041 14603
rect 24075 14600 24087 14603
rect 25682 14600 25688 14612
rect 24075 14572 25688 14600
rect 24075 14569 24087 14572
rect 24029 14563 24087 14569
rect 25682 14560 25688 14572
rect 25740 14560 25746 14612
rect 27154 14560 27160 14612
rect 27212 14560 27218 14612
rect 24854 14492 24860 14544
rect 24912 14532 24918 14544
rect 26326 14532 26332 14544
rect 24912 14504 26332 14532
rect 24912 14492 24918 14504
rect 26326 14492 26332 14504
rect 26384 14492 26390 14544
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19392 14436 19993 14464
rect 19392 14424 19398 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 20220 14436 21189 14464
rect 20220 14424 20226 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22152 14436 22293 14464
rect 22152 14424 22158 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 19889 14399 19947 14405
rect 19889 14396 19901 14399
rect 18984 14368 19901 14396
rect 16853 14359 16911 14365
rect 19889 14365 19901 14368
rect 19935 14396 19947 14399
rect 21358 14396 21364 14408
rect 19935 14368 21364 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 4154 14288 4160 14340
rect 4212 14328 4218 14340
rect 5368 14328 5396 14356
rect 4212 14300 5396 14328
rect 4212 14288 4218 14300
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 5592 14300 6118 14328
rect 5592 14288 5598 14300
rect 7742 14288 7748 14340
rect 7800 14328 7806 14340
rect 12253 14331 12311 14337
rect 7800 14300 12204 14328
rect 7800 14288 7806 14300
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3384 14232 3801 14260
rect 3384 14220 3390 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4430 14220 4436 14272
rect 4488 14260 4494 14272
rect 4525 14263 4583 14269
rect 4525 14260 4537 14263
rect 4488 14232 4537 14260
rect 4488 14220 4494 14232
rect 4525 14229 4537 14232
rect 4571 14229 4583 14263
rect 4525 14223 4583 14229
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 4798 14260 4804 14272
rect 4663 14232 4804 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7837 14263 7895 14269
rect 7837 14260 7849 14263
rect 7340 14232 7849 14260
rect 7340 14220 7346 14232
rect 7837 14229 7849 14232
rect 7883 14229 7895 14263
rect 7837 14223 7895 14229
rect 8205 14263 8263 14269
rect 8205 14229 8217 14263
rect 8251 14260 8263 14263
rect 8478 14260 8484 14272
rect 8251 14232 8484 14260
rect 8251 14229 8263 14232
rect 8205 14223 8263 14229
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8904 14232 9045 14260
rect 8904 14220 8910 14232
rect 9033 14229 9045 14232
rect 9079 14260 9091 14263
rect 9582 14260 9588 14272
rect 9079 14232 9588 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 9916 14232 10609 14260
rect 9916 14220 9922 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 10965 14263 11023 14269
rect 10965 14229 10977 14263
rect 11011 14260 11023 14263
rect 11054 14260 11060 14272
rect 11011 14232 11060 14260
rect 11011 14229 11023 14232
rect 10965 14223 11023 14229
rect 11054 14220 11060 14232
rect 11112 14260 11118 14272
rect 11698 14260 11704 14272
rect 11112 14232 11704 14260
rect 11112 14220 11118 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12176 14260 12204 14300
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 12526 14328 12532 14340
rect 12299 14300 12532 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 13722 14328 13728 14340
rect 13478 14300 13728 14328
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 16298 14328 16304 14340
rect 16146 14300 16304 14328
rect 16298 14288 16304 14300
rect 16356 14288 16362 14340
rect 15930 14260 15936 14272
rect 12176 14232 15936 14260
rect 15930 14220 15936 14232
rect 15988 14260 15994 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15988 14232 16405 14260
rect 15988 14220 15994 14232
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16868 14260 16896 14359
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 23658 14356 23664 14408
rect 23716 14356 23722 14408
rect 23934 14356 23940 14408
rect 23992 14396 23998 14408
rect 26513 14399 26571 14405
rect 26513 14396 26525 14399
rect 23992 14368 26525 14396
rect 23992 14356 23998 14368
rect 26513 14365 26525 14368
rect 26559 14365 26571 14399
rect 26513 14359 26571 14365
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 17092 14300 17618 14328
rect 17092 14288 17098 14300
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 18748 14300 20668 14328
rect 18748 14288 18754 14300
rect 17126 14260 17132 14272
rect 16868 14232 17132 14260
rect 16393 14223 16451 14229
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 19058 14220 19064 14272
rect 19116 14260 19122 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19116 14232 19441 14260
rect 19116 14220 19122 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 19797 14263 19855 14269
rect 19797 14229 19809 14263
rect 19843 14260 19855 14263
rect 19978 14260 19984 14272
rect 19843 14232 19984 14260
rect 19843 14229 19855 14232
rect 19797 14223 19855 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20640 14269 20668 14300
rect 20990 14288 20996 14340
rect 21048 14288 21054 14340
rect 21174 14288 21180 14340
rect 21232 14328 21238 14340
rect 21729 14331 21787 14337
rect 21729 14328 21741 14331
rect 21232 14300 21741 14328
rect 21232 14288 21238 14300
rect 21729 14297 21741 14300
rect 21775 14297 21787 14331
rect 21729 14291 21787 14297
rect 21818 14288 21824 14340
rect 21876 14328 21882 14340
rect 22462 14328 22468 14340
rect 21876 14300 22468 14328
rect 21876 14288 21882 14300
rect 22462 14288 22468 14300
rect 22520 14288 22526 14340
rect 22554 14288 22560 14340
rect 22612 14288 22618 14340
rect 24857 14331 24915 14337
rect 24857 14328 24869 14331
rect 23860 14300 24869 14328
rect 20625 14263 20683 14269
rect 20625 14229 20637 14263
rect 20671 14229 20683 14263
rect 20625 14223 20683 14229
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20956 14232 21097 14260
rect 20956 14220 20962 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 22480 14260 22508 14288
rect 23860 14260 23888 14300
rect 24857 14297 24869 14300
rect 24903 14328 24915 14331
rect 25133 14331 25191 14337
rect 25133 14328 25145 14331
rect 24903 14300 25145 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 25133 14297 25145 14300
rect 25179 14297 25191 14331
rect 25133 14291 25191 14297
rect 25958 14288 25964 14340
rect 26016 14288 26022 14340
rect 22480 14232 23888 14260
rect 21085 14223 21143 14229
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 24673 14263 24731 14269
rect 24673 14229 24685 14263
rect 24719 14260 24731 14263
rect 24946 14260 24952 14272
rect 24719 14232 24952 14260
rect 24719 14229 24731 14232
rect 24673 14223 24731 14229
rect 24946 14220 24952 14232
rect 25004 14260 25010 14272
rect 26510 14260 26516 14272
rect 25004 14232 26516 14260
rect 25004 14220 25010 14232
rect 26510 14220 26516 14232
rect 26568 14220 26574 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3510 14016 3516 14068
rect 3568 14016 3574 14068
rect 5810 14056 5816 14068
rect 3712 14028 5816 14056
rect 106 13880 112 13932
rect 164 13920 170 13932
rect 750 13920 756 13932
rect 164 13892 756 13920
rect 164 13880 170 13892
rect 750 13880 756 13892
rect 808 13880 814 13932
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 3602 13920 3608 13932
rect 1811 13892 3608 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 3712 13929 3740 14028
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6454 14016 6460 14068
rect 6512 14016 6518 14068
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 7892 14028 8125 14056
rect 7892 14016 7898 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 8113 14019 8171 14025
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 8352 14028 8493 14056
rect 8352 14016 8358 14028
rect 8481 14025 8493 14028
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 8570 14016 8576 14068
rect 8628 14016 8634 14068
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 10226 14056 10232 14068
rect 8996 14028 10232 14056
rect 8996 14016 9002 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10376 14028 11069 14056
rect 10376 14016 10382 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12894 14056 12900 14068
rect 11664 14028 12900 14056
rect 11664 14016 11670 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 13262 14056 13268 14068
rect 13127 14028 13268 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 13412 14028 14565 14056
rect 13412 14016 13418 14028
rect 14553 14025 14565 14028
rect 14599 14025 14611 14059
rect 14553 14019 14611 14025
rect 15286 14016 15292 14068
rect 15344 14056 15350 14068
rect 15381 14059 15439 14065
rect 15381 14056 15393 14059
rect 15344 14028 15393 14056
rect 15344 14016 15350 14028
rect 15381 14025 15393 14028
rect 15427 14025 15439 14059
rect 15381 14019 15439 14025
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16390 14056 16396 14068
rect 15887 14028 16396 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17276 14028 18736 14056
rect 17276 14016 17282 14028
rect 5074 13948 5080 14000
rect 5132 13948 5138 14000
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4982 13852 4988 13864
rect 4479 13824 4988 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5552 13852 5580 13880
rect 5132 13824 5580 13852
rect 5132 13812 5138 13824
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 5905 13855 5963 13861
rect 5905 13852 5917 13855
rect 5684 13824 5917 13852
rect 5684 13812 5690 13824
rect 5905 13821 5917 13824
rect 5951 13852 5963 13855
rect 6178 13852 6184 13864
rect 5951 13824 6184 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6472 13852 6500 14016
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 6696 13960 7389 13988
rect 6696 13948 6702 13960
rect 7377 13957 7389 13960
rect 7423 13957 7435 13991
rect 7377 13951 7435 13957
rect 8754 13948 8760 14000
rect 8812 13988 8818 14000
rect 9490 13988 9496 14000
rect 8812 13960 9496 13988
rect 8812 13948 8818 13960
rect 9490 13948 9496 13960
rect 9548 13988 9554 14000
rect 13538 13988 13544 14000
rect 9548 13960 10074 13988
rect 11716 13960 13544 13988
rect 9548 13948 9554 13960
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 11716 13929 11744 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 13872 13960 15761 13988
rect 13872 13948 13878 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 16761 13991 16819 13997
rect 16761 13988 16773 13991
rect 16356 13960 16773 13988
rect 16356 13948 16362 13960
rect 16761 13957 16773 13960
rect 16807 13988 16819 13991
rect 17034 13988 17040 14000
rect 16807 13960 17040 13988
rect 16807 13957 16819 13960
rect 16761 13951 16819 13957
rect 17034 13948 17040 13960
rect 17092 13988 17098 14000
rect 17862 13988 17868 14000
rect 17092 13960 17868 13988
rect 17092 13948 17098 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 18708 13988 18736 14028
rect 18874 14016 18880 14068
rect 18932 14016 18938 14068
rect 19242 14016 19248 14068
rect 19300 14016 19306 14068
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 20438 14056 20444 14068
rect 19567 14028 20444 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 20622 14016 20628 14068
rect 20680 14016 20686 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 21048 14028 21373 14056
rect 21048 14016 21054 14028
rect 21361 14025 21373 14028
rect 21407 14056 21419 14059
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 21407 14028 21557 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21545 14025 21557 14028
rect 21591 14056 21603 14059
rect 22462 14056 22468 14068
rect 21591 14028 22468 14056
rect 21591 14025 21603 14028
rect 21545 14019 21603 14025
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14025 23259 14059
rect 23201 14019 23259 14025
rect 20640 13988 20668 14016
rect 18708 13960 20668 13988
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 23216 13988 23244 14019
rect 24118 14016 24124 14068
rect 24176 14056 24182 14068
rect 24397 14059 24455 14065
rect 24397 14056 24409 14059
rect 24176 14028 24409 14056
rect 24176 14016 24182 14028
rect 24397 14025 24409 14028
rect 24443 14025 24455 14059
rect 24397 14019 24455 14025
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 26142 14056 26148 14068
rect 25556 14028 26148 14056
rect 25556 14016 25562 14028
rect 26142 14016 26148 14028
rect 26200 14056 26206 14068
rect 26237 14059 26295 14065
rect 26237 14056 26249 14059
rect 26200 14028 26249 14056
rect 26200 14016 26206 14028
rect 26237 14025 26249 14028
rect 26283 14025 26295 14059
rect 26237 14019 26295 14025
rect 26326 14016 26332 14068
rect 26384 14056 26390 14068
rect 26697 14059 26755 14065
rect 26697 14056 26709 14059
rect 26384 14028 26709 14056
rect 26384 14016 26390 14028
rect 26697 14025 26709 14028
rect 26743 14056 26755 14059
rect 27706 14056 27712 14068
rect 26743 14028 27712 14056
rect 26743 14025 26755 14028
rect 26697 14019 26755 14025
rect 27706 14016 27712 14028
rect 27764 14016 27770 14068
rect 20772 13960 23244 13988
rect 23661 13991 23719 13997
rect 20772 13948 20778 13960
rect 23661 13957 23673 13991
rect 23707 13988 23719 13991
rect 24854 13988 24860 14000
rect 23707 13960 24860 13988
rect 23707 13957 23719 13960
rect 23661 13951 23719 13957
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 25409 13991 25467 13997
rect 25409 13957 25421 13991
rect 25455 13988 25467 13991
rect 25590 13988 25596 14000
rect 25455 13960 25596 13988
rect 25455 13957 25467 13960
rect 25409 13951 25467 13957
rect 25590 13948 25596 13960
rect 25648 13988 25654 14000
rect 26053 13991 26111 13997
rect 26053 13988 26065 13991
rect 25648 13960 26065 13988
rect 25648 13948 25654 13960
rect 26053 13957 26065 13960
rect 26099 13957 26111 13991
rect 26053 13951 26111 13957
rect 11701 13923 11759 13929
rect 7800 13892 9260 13920
rect 7800 13880 7806 13892
rect 6420 13824 6500 13852
rect 6420 13812 6426 13824
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 6822 13852 6828 13864
rect 6696 13824 6828 13852
rect 6696 13812 6702 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7558 13812 7564 13864
rect 7616 13812 7622 13864
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 750 13744 756 13796
rect 808 13784 814 13796
rect 1210 13784 1216 13796
rect 808 13756 1216 13784
rect 808 13744 814 13756
rect 1210 13744 1216 13756
rect 1268 13744 1274 13796
rect 8478 13784 8484 13796
rect 5460 13756 8484 13784
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 5460 13716 5488 13756
rect 8478 13744 8484 13756
rect 8536 13744 8542 13796
rect 8772 13784 8800 13815
rect 9232 13784 9260 13892
rect 11701 13889 11713 13923
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12158 13920 12164 13932
rect 12023 13892 12164 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 15654 13920 15660 13932
rect 14507 13892 15660 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 20530 13880 20536 13932
rect 20588 13880 20594 13932
rect 20625 13923 20683 13929
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 20671 13892 22094 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9582 13852 9588 13864
rect 9416 13824 9588 13852
rect 9416 13784 9444 13824
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10284 13824 12664 13852
rect 10284 13812 10290 13824
rect 8772 13756 8892 13784
rect 9232 13756 9444 13784
rect 3844 13688 5488 13716
rect 3844 13676 3850 13688
rect 6914 13676 6920 13728
rect 6972 13676 6978 13728
rect 8864 13716 8892 13756
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 12342 13784 12348 13796
rect 11020 13756 12348 13784
rect 11020 13744 11026 13756
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 9582 13716 9588 13728
rect 8864 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13716 9646 13728
rect 10318 13716 10324 13728
rect 9640 13688 10324 13716
rect 9640 13676 9646 13688
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 12636 13716 12664 13824
rect 12894 13812 12900 13864
rect 12952 13812 12958 13864
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13311 13824 13553 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13541 13821 13553 13824
rect 13587 13852 13599 13855
rect 13722 13852 13728 13864
rect 13587 13824 13728 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 15378 13852 15384 13864
rect 14783 13824 15384 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15930 13812 15936 13864
rect 15988 13812 15994 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17236 13824 17417 13852
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13814 13784 13820 13796
rect 12768 13756 13820 13784
rect 12768 13744 12774 13756
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13784 14151 13787
rect 14366 13784 14372 13796
rect 14139 13756 14372 13784
rect 14139 13753 14151 13756
rect 14093 13747 14151 13753
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 16482 13744 16488 13796
rect 16540 13784 16546 13796
rect 17236 13784 17264 13824
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 17494 13812 17500 13864
rect 17552 13852 17558 13864
rect 20809 13855 20867 13861
rect 17552 13824 20208 13852
rect 17552 13812 17558 13824
rect 16540 13756 17264 13784
rect 16540 13744 16546 13756
rect 18506 13744 18512 13796
rect 18564 13784 18570 13796
rect 18966 13784 18972 13796
rect 18564 13756 18972 13784
rect 18564 13744 18570 13756
rect 18966 13744 18972 13756
rect 19024 13744 19030 13796
rect 20180 13793 20208 13824
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13753 20223 13787
rect 20824 13784 20852 13815
rect 20898 13812 20904 13864
rect 20956 13852 20962 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 20956 13824 21189 13852
rect 20956 13812 20962 13824
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 22066 13852 22094 13892
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22244 13892 22385 13920
rect 22244 13880 22250 13892
rect 22373 13889 22385 13892
rect 22419 13889 22431 13923
rect 23474 13920 23480 13932
rect 22373 13883 22431 13889
rect 22480 13892 23480 13920
rect 22480 13852 22508 13892
rect 23474 13880 23480 13892
rect 23532 13880 23538 13932
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13920 23627 13923
rect 23615 13892 24348 13920
rect 23615 13889 23627 13892
rect 23569 13883 23627 13889
rect 24320 13864 24348 13892
rect 24578 13880 24584 13932
rect 24636 13880 24642 13932
rect 26513 13923 26571 13929
rect 26513 13920 26525 13923
rect 24688 13892 26525 13920
rect 22066 13824 22508 13852
rect 22557 13855 22615 13861
rect 21177 13815 21235 13821
rect 22557 13821 22569 13855
rect 22603 13821 22615 13855
rect 22557 13815 22615 13821
rect 23753 13855 23811 13861
rect 23753 13821 23765 13855
rect 23799 13821 23811 13855
rect 23753 13815 23811 13821
rect 21818 13784 21824 13796
rect 20824 13756 21824 13784
rect 20165 13747 20223 13753
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 22572 13784 22600 13815
rect 22646 13784 22652 13796
rect 22572 13756 22652 13784
rect 22646 13744 22652 13756
rect 22704 13784 22710 13796
rect 23768 13784 23796 13815
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24688 13852 24716 13892
rect 26513 13889 26525 13892
rect 26559 13920 26571 13923
rect 30374 13920 30380 13932
rect 26559 13892 30380 13920
rect 26559 13889 26571 13892
rect 26513 13883 26571 13889
rect 30374 13880 30380 13892
rect 30432 13880 30438 13932
rect 24360 13824 24716 13852
rect 25685 13855 25743 13861
rect 24360 13812 24366 13824
rect 25685 13821 25697 13855
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 22704 13756 23796 13784
rect 22704 13744 22710 13756
rect 24486 13744 24492 13796
rect 24544 13784 24550 13796
rect 24946 13784 24952 13796
rect 24544 13756 24952 13784
rect 24544 13744 24550 13756
rect 24946 13744 24952 13756
rect 25004 13744 25010 13796
rect 25700 13784 25728 13815
rect 26234 13784 26240 13796
rect 25700 13756 26240 13784
rect 26234 13744 26240 13756
rect 26292 13744 26298 13796
rect 15654 13716 15660 13728
rect 12636 13688 15660 13716
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 18012 13688 22017 13716
rect 18012 13676 18018 13688
rect 22005 13685 22017 13688
rect 22051 13685 22063 13719
rect 22005 13679 22063 13685
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 23934 13716 23940 13728
rect 22152 13688 23940 13716
rect 22152 13676 22158 13688
rect 23934 13676 23940 13688
rect 23992 13676 23998 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 5994 13512 6000 13524
rect 3651 13484 6000 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 7190 13512 7196 13524
rect 6840 13484 7196 13512
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 3878 13444 3884 13456
rect 3476 13416 3884 13444
rect 3476 13404 3482 13416
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 5074 13444 5080 13456
rect 4479 13416 5080 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 6840 13444 6868 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 14534 13515 14592 13521
rect 14534 13512 14546 13515
rect 7524 13484 14546 13512
rect 7524 13472 7530 13484
rect 14534 13481 14546 13484
rect 14580 13481 14592 13515
rect 14534 13475 14592 13481
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15160 13484 16037 13512
rect 15160 13472 15166 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 20714 13512 20720 13524
rect 17644 13484 20720 13512
rect 17644 13472 17650 13484
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 22005 13515 22063 13521
rect 22005 13481 22017 13515
rect 22051 13512 22063 13515
rect 22094 13512 22100 13524
rect 22051 13484 22100 13512
rect 22051 13481 22063 13484
rect 22005 13475 22063 13481
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22462 13472 22468 13524
rect 22520 13512 22526 13524
rect 22925 13515 22983 13521
rect 22925 13512 22937 13515
rect 22520 13484 22937 13512
rect 22520 13472 22526 13484
rect 22925 13481 22937 13484
rect 22971 13512 22983 13515
rect 23382 13512 23388 13524
rect 22971 13484 23388 13512
rect 22971 13481 22983 13484
rect 22925 13475 22983 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 5316 13416 6868 13444
rect 8573 13447 8631 13453
rect 5316 13404 5322 13416
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 8619 13416 11008 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4893 13379 4951 13385
rect 4893 13376 4905 13379
rect 4672 13348 4905 13376
rect 4672 13336 4678 13348
rect 4893 13345 4905 13348
rect 4939 13345 4951 13379
rect 4893 13339 4951 13345
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5994 13376 6000 13388
rect 5031 13348 6000 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 6178 13336 6184 13388
rect 6236 13336 6242 13388
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7558 13376 7564 13388
rect 7147 13348 7564 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 8588 13376 8616 13407
rect 7800 13348 8616 13376
rect 7800 13336 7806 13348
rect 9766 13336 9772 13388
rect 9824 13336 9830 13388
rect 10980 13385 11008 13416
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 11112 13416 11437 13444
rect 11112 13404 11118 13416
rect 11425 13413 11437 13416
rect 11471 13413 11483 13447
rect 11425 13407 11483 13413
rect 11609 13447 11667 13453
rect 11609 13413 11621 13447
rect 11655 13444 11667 13447
rect 11698 13444 11704 13456
rect 11655 13416 11704 13444
rect 11655 13413 11667 13416
rect 11609 13407 11667 13413
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 13630 13404 13636 13456
rect 13688 13444 13694 13456
rect 13725 13447 13783 13453
rect 13725 13444 13737 13447
rect 13688 13416 13737 13444
rect 13688 13404 13694 13416
rect 13725 13413 13737 13416
rect 13771 13413 13783 13447
rect 13725 13407 13783 13413
rect 15654 13404 15660 13456
rect 15712 13444 15718 13456
rect 16850 13444 16856 13456
rect 15712 13416 16856 13444
rect 15712 13404 15718 13416
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 18877 13447 18935 13453
rect 18877 13444 18889 13447
rect 18656 13416 18889 13444
rect 18656 13404 18662 13416
rect 18877 13413 18889 13416
rect 18923 13413 18935 13447
rect 18877 13407 18935 13413
rect 24302 13404 24308 13456
rect 24360 13444 24366 13456
rect 24581 13447 24639 13453
rect 24581 13444 24593 13447
rect 24360 13416 24593 13444
rect 24360 13404 24366 13416
rect 24581 13413 24593 13416
rect 24627 13413 24639 13447
rect 24581 13407 24639 13413
rect 10965 13379 11023 13385
rect 10704 13348 10916 13376
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 4338 13308 4344 13320
rect 3936 13280 4344 13308
rect 3936 13268 3942 13280
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5442 13308 5448 13320
rect 4847 13280 5448 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5868 13280 6101 13308
rect 5868 13268 5874 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 10704 13308 10732 13348
rect 8536 13280 10732 13308
rect 8536 13268 8542 13280
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10888 13308 10916 13348
rect 10965 13345 10977 13379
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12250 13376 12256 13388
rect 12032 13348 12256 13376
rect 12032 13336 12038 13348
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 12308 13348 14289 13376
rect 12308 13336 12314 13348
rect 14277 13345 14289 13348
rect 14323 13376 14335 13379
rect 14642 13376 14648 13388
rect 14323 13348 14648 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 14642 13336 14648 13348
rect 14700 13376 14706 13388
rect 15102 13376 15108 13388
rect 14700 13348 15108 13376
rect 14700 13336 14706 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 16666 13376 16672 13388
rect 16531 13348 16672 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 19702 13376 19708 13388
rect 17184 13348 19708 13376
rect 17184 13336 17190 13348
rect 19702 13336 19708 13348
rect 19760 13376 19766 13388
rect 20533 13379 20591 13385
rect 19760 13348 20300 13376
rect 19760 13336 19766 13348
rect 20272 13320 20300 13348
rect 20533 13345 20545 13379
rect 20579 13376 20591 13379
rect 20898 13376 20904 13388
rect 20579 13348 20904 13376
rect 20579 13345 20591 13348
rect 20533 13339 20591 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 22186 13336 22192 13388
rect 22244 13376 22250 13388
rect 22244 13348 23704 13376
rect 22244 13336 22250 13348
rect 11330 13308 11336 13320
rect 10888 13280 11336 13308
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 16942 13308 16948 13320
rect 16080 13280 16948 13308
rect 16080 13268 16086 13280
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18472 13280 19901 13308
rect 18472 13268 18478 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 23676 13317 23704 13348
rect 23750 13336 23756 13388
rect 23808 13336 23814 13388
rect 23842 13336 23848 13388
rect 23900 13336 23906 13388
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 23992 13348 25145 13376
rect 23992 13336 23998 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 22649 13311 22707 13317
rect 22649 13308 22661 13311
rect 21968 13280 22661 13308
rect 21968 13268 21974 13280
rect 22649 13277 22661 13280
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13308 23719 13311
rect 24394 13308 24400 13320
rect 23707 13280 24400 13308
rect 23707 13277 23719 13280
rect 23661 13271 23719 13277
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25038 13308 25044 13320
rect 24995 13280 25044 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 25777 13311 25835 13317
rect 25777 13308 25789 13311
rect 25740 13280 25789 13308
rect 25740 13268 25746 13280
rect 25777 13277 25789 13280
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 3973 13243 4031 13249
rect 3973 13209 3985 13243
rect 4019 13240 4031 13243
rect 6270 13240 6276 13252
rect 4019 13212 6276 13240
rect 4019 13209 4031 13212
rect 3973 13203 4031 13209
rect 6270 13200 6276 13212
rect 6328 13200 6334 13252
rect 7190 13200 7196 13252
rect 7248 13240 7254 13252
rect 10689 13243 10747 13249
rect 7248 13212 7590 13240
rect 7248 13200 7254 13212
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 10735 13212 11652 13240
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4430 13172 4436 13184
rect 4203 13144 4436 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5718 13172 5724 13184
rect 5675 13144 5724 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 5868 13144 6009 13172
rect 5868 13132 5874 13144
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9214 13172 9220 13184
rect 9171 13144 9220 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9585 13175 9643 13181
rect 9585 13141 9597 13175
rect 9631 13172 9643 13175
rect 10134 13172 10140 13184
rect 9631 13144 10140 13172
rect 9631 13141 9643 13144
rect 9585 13135 9643 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 10318 13132 10324 13184
rect 10376 13132 10382 13184
rect 11624 13172 11652 13212
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12253 13243 12311 13249
rect 12253 13240 12265 13243
rect 11756 13212 12265 13240
rect 11756 13200 11762 13212
rect 12253 13209 12265 13212
rect 12299 13209 12311 13243
rect 13722 13240 13728 13252
rect 13478 13212 13728 13240
rect 12253 13203 12311 13209
rect 13722 13200 13728 13212
rect 13780 13240 13786 13252
rect 16666 13240 16672 13252
rect 13780 13212 15042 13240
rect 15856 13212 16672 13240
rect 13780 13200 13786 13212
rect 13998 13172 14004 13184
rect 11624 13144 14004 13172
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14936 13172 14964 13212
rect 15856 13172 15884 13212
rect 16666 13200 16672 13212
rect 16724 13200 16730 13252
rect 17405 13243 17463 13249
rect 17405 13209 17417 13243
rect 17451 13240 17463 13243
rect 17451 13212 17816 13240
rect 17451 13209 17463 13212
rect 17405 13203 17463 13209
rect 17788 13184 17816 13212
rect 18046 13200 18052 13252
rect 18104 13200 18110 13252
rect 21082 13200 21088 13252
rect 21140 13200 21146 13252
rect 32214 13240 32220 13252
rect 22480 13212 32220 13240
rect 14936 13144 15884 13172
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 17310 13172 17316 13184
rect 15988 13144 17316 13172
rect 15988 13132 15994 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 17770 13132 17776 13184
rect 17828 13132 17834 13184
rect 18322 13132 18328 13184
rect 18380 13172 18386 13184
rect 22480 13181 22508 13212
rect 32214 13200 32220 13212
rect 32272 13200 32278 13252
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 18380 13144 19441 13172
rect 18380 13132 18386 13144
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 22465 13175 22523 13181
rect 22465 13141 22477 13175
rect 22511 13141 22523 13175
rect 22465 13135 22523 13141
rect 23290 13132 23296 13184
rect 23348 13132 23354 13184
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 24486 13172 24492 13184
rect 23716 13144 24492 13172
rect 23716 13132 23722 13144
rect 24486 13132 24492 13144
rect 24544 13132 24550 13184
rect 25041 13175 25099 13181
rect 25041 13141 25053 13175
rect 25087 13172 25099 13175
rect 25774 13172 25780 13184
rect 25087 13144 25780 13172
rect 25087 13141 25099 13144
rect 25041 13135 25099 13141
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 26418 13132 26424 13184
rect 26476 13132 26482 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 3326 12968 3332 12980
rect 2915 12940 3332 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3326 12928 3332 12940
rect 3384 12968 3390 12980
rect 3384 12940 4200 12968
rect 3384 12928 3390 12940
rect 3786 12860 3792 12912
rect 3844 12860 3850 12912
rect 4172 12900 4200 12940
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 5534 12968 5540 12980
rect 5408 12940 5540 12968
rect 5408 12928 5414 12940
rect 5534 12928 5540 12940
rect 5592 12968 5598 12980
rect 5592 12940 6868 12968
rect 5592 12928 5598 12940
rect 6840 12912 6868 12940
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7285 12971 7343 12977
rect 7285 12968 7297 12971
rect 6972 12940 7297 12968
rect 6972 12928 6978 12940
rect 7285 12937 7297 12940
rect 7331 12937 7343 12971
rect 9306 12968 9312 12980
rect 7285 12931 7343 12937
rect 8128 12940 9312 12968
rect 4982 12900 4988 12912
rect 4172 12872 4988 12900
rect 4982 12860 4988 12872
rect 5040 12860 5046 12912
rect 6086 12860 6092 12912
rect 6144 12900 6150 12912
rect 6365 12903 6423 12909
rect 6365 12900 6377 12903
rect 6144 12872 6377 12900
rect 6144 12860 6150 12872
rect 6365 12869 6377 12872
rect 6411 12869 6423 12903
rect 6365 12863 6423 12869
rect 6822 12860 6828 12912
rect 6880 12900 6886 12912
rect 8128 12900 8156 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 10652 12940 11008 12968
rect 10652 12928 10658 12940
rect 6880 12872 8156 12900
rect 6880 12860 6886 12872
rect 1118 12792 1124 12844
rect 1176 12832 1182 12844
rect 1486 12832 1492 12844
rect 1176 12804 1492 12832
rect 1176 12792 1182 12804
rect 1486 12792 1492 12804
rect 1544 12832 1550 12844
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 1544 12804 1593 12832
rect 1544 12792 1550 12804
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12832 3203 12835
rect 3602 12832 3608 12844
rect 3191 12804 3608 12832
rect 3191 12801 3203 12804
rect 3145 12795 3203 12801
rect 3602 12792 3608 12804
rect 3660 12792 3666 12844
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4249 12835 4307 12841
rect 4249 12832 4261 12835
rect 4120 12804 4261 12832
rect 4120 12792 4126 12804
rect 4249 12801 4261 12804
rect 4295 12801 4307 12835
rect 6178 12832 6184 12844
rect 4249 12795 4307 12801
rect 5828 12804 6184 12832
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12733 1915 12767
rect 1857 12727 1915 12733
rect 1872 12628 1900 12727
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 4154 12764 4160 12776
rect 2740 12736 4160 12764
rect 2740 12724 2746 12736
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5828 12764 5856 12804
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6788 12804 7389 12832
rect 6788 12792 6794 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7742 12832 7748 12844
rect 7377 12795 7435 12801
rect 7576 12804 7748 12832
rect 4571 12736 5856 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5994 12724 6000 12776
rect 6052 12724 6058 12776
rect 7576 12773 7604 12804
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 8128 12841 8156 12872
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12900 10195 12903
rect 10410 12900 10416 12912
rect 10183 12872 10416 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 10870 12900 10876 12912
rect 10560 12872 10876 12900
rect 10560 12860 10566 12872
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10284 12804 10609 12832
rect 10284 12792 10290 12804
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 10980 12832 11008 12940
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 12768 12940 12817 12968
rect 12768 12928 12774 12940
rect 12805 12937 12817 12940
rect 12851 12937 12863 12971
rect 12805 12931 12863 12937
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 15194 12968 15200 12980
rect 14415 12940 15200 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 15562 12928 15568 12980
rect 15620 12928 15626 12980
rect 16025 12971 16083 12977
rect 16025 12937 16037 12971
rect 16071 12968 16083 12971
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16071 12940 17141 12968
rect 16071 12937 16083 12940
rect 16025 12931 16083 12937
rect 17129 12937 17141 12940
rect 17175 12937 17187 12971
rect 17129 12931 17187 12937
rect 17494 12928 17500 12980
rect 17552 12928 17558 12980
rect 17586 12928 17592 12980
rect 17644 12928 17650 12980
rect 18693 12971 18751 12977
rect 18693 12937 18705 12971
rect 18739 12968 18751 12971
rect 23290 12968 23296 12980
rect 18739 12940 23296 12968
rect 18739 12937 18751 12940
rect 18693 12931 18751 12937
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 14737 12903 14795 12909
rect 13004 12872 14136 12900
rect 13004 12832 13032 12872
rect 10827 12804 13032 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 14108 12841 14136 12872
rect 14737 12869 14749 12903
rect 14783 12900 14795 12903
rect 14783 12872 18644 12900
rect 14783 12869 14795 12872
rect 14737 12863 14795 12869
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13412 12804 13461 12832
rect 13412 12792 13418 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 14139 12804 14872 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 7561 12767 7619 12773
rect 7561 12764 7573 12767
rect 6748 12736 7573 12764
rect 6748 12708 6776 12736
rect 7561 12733 7573 12736
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 7708 12736 8401 12764
rect 7708 12724 7714 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 9508 12764 9536 12792
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 9508 12736 10977 12764
rect 6730 12656 6736 12708
rect 6788 12656 6794 12708
rect 6917 12699 6975 12705
rect 6917 12665 6929 12699
rect 6963 12696 6975 12699
rect 6963 12668 7052 12696
rect 6963 12665 6975 12668
rect 6917 12659 6975 12665
rect 6546 12628 6552 12640
rect 1872 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7024 12628 7052 12668
rect 7742 12628 7748 12640
rect 7024 12600 7748 12628
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 9508 12628 9536 12736
rect 10965 12733 10977 12736
rect 11011 12764 11023 12767
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11011 12736 11253 12764
rect 11011 12733 11023 12736
rect 10965 12727 11023 12733
rect 11241 12733 11253 12736
rect 11287 12733 11299 12767
rect 12802 12764 12808 12776
rect 11241 12727 11299 12733
rect 12084 12736 12808 12764
rect 11517 12699 11575 12705
rect 11517 12696 11529 12699
rect 10980 12668 11529 12696
rect 10980 12640 11008 12668
rect 11517 12665 11529 12668
rect 11563 12665 11575 12699
rect 11517 12659 11575 12665
rect 8444 12600 9536 12628
rect 8444 12588 8450 12600
rect 10962 12588 10968 12640
rect 11020 12588 11026 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 12084 12637 12112 12736
rect 12802 12724 12808 12736
rect 12860 12764 12866 12776
rect 14844 12773 14872 12804
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15528 12804 15945 12832
rect 15528 12792 15534 12804
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 18506 12832 18512 12844
rect 15933 12795 15991 12801
rect 16132 12804 18512 12832
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12860 12736 12909 12764
rect 12860 12724 12866 12736
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 14918 12764 14924 12776
rect 14875 12736 14924 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 12342 12656 12348 12708
rect 12400 12696 12406 12708
rect 13096 12696 13124 12727
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 16132 12764 16160 12804
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 18616 12832 18644 12872
rect 19518 12860 19524 12912
rect 19576 12860 19582 12912
rect 20254 12860 20260 12912
rect 20312 12860 20318 12912
rect 20714 12860 20720 12912
rect 20772 12900 20778 12912
rect 20901 12903 20959 12909
rect 20901 12900 20913 12903
rect 20772 12872 20913 12900
rect 20772 12860 20778 12872
rect 20901 12869 20913 12872
rect 20947 12869 20959 12903
rect 20901 12863 20959 12869
rect 21637 12903 21695 12909
rect 21637 12869 21649 12903
rect 21683 12900 21695 12903
rect 22186 12900 22192 12912
rect 21683 12872 22192 12900
rect 21683 12869 21695 12872
rect 21637 12863 21695 12869
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 23198 12900 23204 12912
rect 22664 12872 23204 12900
rect 18616 12804 19104 12832
rect 15059 12736 16160 12764
rect 16209 12767 16267 12773
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 16209 12733 16221 12767
rect 16255 12764 16267 12767
rect 16255 12736 16620 12764
rect 16255 12733 16267 12736
rect 16209 12727 16267 12733
rect 15930 12696 15936 12708
rect 12400 12668 15936 12696
rect 12400 12656 12406 12668
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11388 12600 12081 12628
rect 11388 12588 11394 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 12710 12628 12716 12640
rect 12483 12600 12716 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 13817 12631 13875 12637
rect 13817 12628 13829 12631
rect 13780 12600 13829 12628
rect 13780 12588 13786 12600
rect 13817 12597 13829 12600
rect 13863 12628 13875 12631
rect 14366 12628 14372 12640
rect 13863 12600 14372 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 16592 12628 16620 12736
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 17034 12764 17040 12776
rect 16724 12736 17040 12764
rect 16724 12724 16730 12736
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 17681 12767 17739 12773
rect 17681 12764 17693 12767
rect 17644 12736 17693 12764
rect 17644 12724 17650 12736
rect 17681 12733 17693 12736
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 18785 12767 18843 12773
rect 18785 12733 18797 12767
rect 18831 12764 18843 12767
rect 18831 12736 18920 12764
rect 18831 12733 18843 12736
rect 18785 12727 18843 12733
rect 18230 12628 18236 12640
rect 16592 12600 18236 12628
rect 18230 12588 18236 12600
rect 18288 12588 18294 12640
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 18892 12628 18920 12736
rect 18966 12724 18972 12776
rect 19024 12724 19030 12776
rect 19076 12764 19104 12804
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21450 12832 21456 12844
rect 21140 12804 21456 12832
rect 21140 12792 21146 12804
rect 21450 12792 21456 12804
rect 21508 12832 21514 12844
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 21508 12804 22477 12832
rect 21508 12792 21514 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 22005 12767 22063 12773
rect 22005 12764 22017 12767
rect 19076 12736 22017 12764
rect 22005 12733 22017 12736
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 22664 12628 22692 12872
rect 23198 12860 23204 12872
rect 23256 12860 23262 12912
rect 23750 12860 23756 12912
rect 23808 12860 23814 12912
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12832 25283 12835
rect 26234 12832 26240 12844
rect 25271 12804 26240 12832
rect 25271 12801 25283 12804
rect 25225 12795 25283 12801
rect 26234 12792 26240 12804
rect 26292 12792 26298 12844
rect 23017 12767 23075 12773
rect 23017 12733 23029 12767
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 26418 12764 26424 12776
rect 23339 12736 26424 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 18892 12600 22692 12628
rect 23032 12628 23060 12727
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 23382 12628 23388 12640
rect 23032 12600 23388 12628
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 24670 12588 24676 12640
rect 24728 12628 24734 12640
rect 24765 12631 24823 12637
rect 24765 12628 24777 12631
rect 24728 12600 24777 12628
rect 24728 12588 24734 12600
rect 24765 12597 24777 12600
rect 24811 12597 24823 12631
rect 24765 12591 24823 12597
rect 25866 12588 25872 12640
rect 25924 12588 25930 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 2406 12424 2412 12436
rect 2363 12396 2412 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4062 12424 4068 12436
rect 3660 12396 4068 12424
rect 3660 12384 3666 12396
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4157 12427 4215 12433
rect 4157 12393 4169 12427
rect 4203 12424 4215 12427
rect 4890 12424 4896 12436
rect 4203 12396 4896 12424
rect 4203 12393 4215 12396
rect 4157 12387 4215 12393
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5077 12427 5135 12433
rect 5077 12393 5089 12427
rect 5123 12424 5135 12427
rect 7650 12424 7656 12436
rect 5123 12396 7656 12424
rect 5123 12393 5135 12396
rect 5077 12387 5135 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 10870 12424 10876 12436
rect 8312 12396 10876 12424
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 3476 12328 5672 12356
rect 3476 12316 3482 12328
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 5442 12288 5448 12300
rect 3844 12260 5448 12288
rect 3844 12248 3850 12260
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5534 12248 5540 12300
rect 5592 12248 5598 12300
rect 5644 12288 5672 12328
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 8312 12356 8340 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 11020 12396 14473 12424
rect 11020 12384 11026 12396
rect 14461 12393 14473 12396
rect 14507 12424 14519 12427
rect 14734 12424 14740 12436
rect 14507 12396 14740 12424
rect 14507 12393 14519 12396
rect 14461 12387 14519 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 15436 12396 17969 12424
rect 15436 12384 15442 12396
rect 17957 12393 17969 12396
rect 18003 12424 18015 12427
rect 18230 12424 18236 12436
rect 18003 12396 18236 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 18230 12384 18236 12396
rect 18288 12424 18294 12436
rect 18782 12424 18788 12436
rect 18288 12396 18788 12424
rect 18288 12384 18294 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19444 12396 22094 12424
rect 12066 12356 12072 12368
rect 7248 12328 8340 12356
rect 8404 12328 12072 12356
rect 7248 12316 7254 12328
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5644 12260 5825 12288
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 6420 12260 7512 12288
rect 6420 12248 6426 12260
rect 1670 12180 1676 12232
rect 1728 12180 1734 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 3142 12220 3148 12232
rect 2823 12192 3148 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 3421 12223 3479 12229
rect 3421 12220 3433 12223
rect 3292 12192 3433 12220
rect 3292 12180 3298 12192
rect 3421 12189 3433 12192
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 7484 12220 7512 12260
rect 7558 12248 7564 12300
rect 7616 12248 7622 12300
rect 8404 12297 8432 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 13998 12356 14004 12368
rect 12452 12328 14004 12356
rect 8389 12291 8447 12297
rect 8389 12257 8401 12291
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9364 12260 9873 12288
rect 9364 12248 9370 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 12452 12297 12480 12328
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 14090 12316 14096 12368
rect 14148 12316 14154 12368
rect 17494 12316 17500 12368
rect 17552 12356 17558 12368
rect 18601 12359 18659 12365
rect 18601 12356 18613 12359
rect 17552 12328 18613 12356
rect 17552 12316 17558 12328
rect 18601 12325 18613 12328
rect 18647 12325 18659 12359
rect 19058 12356 19064 12368
rect 18601 12319 18659 12325
rect 18708 12328 19064 12356
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10928 12260 11161 12288
rect 10928 12248 10934 12260
rect 11149 12257 11161 12260
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13679 12260 14504 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 8938 12220 8944 12232
rect 4479 12192 5580 12220
rect 7484 12192 8944 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 5552 12152 5580 12192
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 10284 12192 12173 12220
rect 10284 12180 10290 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14476 12220 14504 12260
rect 14660 12260 15148 12288
rect 14660 12220 14688 12260
rect 13495 12192 14412 12220
rect 14476 12192 14688 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 2004 12124 5212 12152
rect 5552 12124 6224 12152
rect 2004 12112 2010 12124
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 4338 12084 4344 12096
rect 4019 12056 4344 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 4338 12044 4344 12056
rect 4396 12084 4402 12096
rect 4982 12084 4988 12096
rect 4396 12056 4988 12084
rect 4396 12044 4402 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5184 12084 5212 12124
rect 5994 12084 6000 12096
rect 5184 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6196 12084 6224 12124
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 7374 12112 7380 12164
rect 7432 12152 7438 12164
rect 7432 12124 7604 12152
rect 7432 12112 7438 12124
rect 7466 12084 7472 12096
rect 6196 12056 7472 12084
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7576 12084 7604 12124
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 7708 12124 8524 12152
rect 7708 12112 7714 12124
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7576 12056 7849 12084
rect 7837 12053 7849 12056
rect 7883 12084 7895 12087
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7883 12056 8033 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 8021 12053 8033 12056
rect 8067 12084 8079 12087
rect 8386 12084 8392 12096
rect 8067 12056 8392 12084
rect 8067 12053 8079 12056
rect 8021 12047 8079 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8496 12084 8524 12124
rect 10410 12112 10416 12164
rect 10468 12152 10474 12164
rect 11057 12155 11115 12161
rect 11057 12152 11069 12155
rect 10468 12124 11069 12152
rect 10468 12112 10474 12124
rect 11057 12121 11069 12124
rect 11103 12121 11115 12155
rect 11057 12115 11115 12121
rect 12253 12155 12311 12161
rect 12253 12121 12265 12155
rect 12299 12152 12311 12155
rect 13814 12152 13820 12164
rect 12299 12124 13820 12152
rect 12299 12121 12311 12124
rect 12253 12115 12311 12121
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 14384 12152 14412 12192
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14792 12192 14841 12220
rect 14792 12180 14798 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 15120 12220 15148 12260
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15565 12291 15623 12297
rect 15565 12288 15577 12291
rect 15252 12260 15577 12288
rect 15252 12248 15258 12260
rect 15565 12257 15577 12260
rect 15611 12288 15623 12291
rect 16209 12291 16267 12297
rect 16209 12288 16221 12291
rect 15611 12260 16221 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 16209 12257 16221 12260
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 18322 12288 18328 12300
rect 17276 12260 18328 12288
rect 17276 12248 17282 12260
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 16114 12220 16120 12232
rect 15120 12192 16120 12220
rect 14829 12183 14887 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 18708 12220 18736 12328
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 19444 12288 19472 12396
rect 22066 12356 22094 12396
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 23290 12424 23296 12436
rect 22796 12396 23296 12424
rect 22796 12384 22802 12396
rect 23290 12384 23296 12396
rect 23348 12424 23354 12436
rect 25958 12424 25964 12436
rect 23348 12396 25964 12424
rect 23348 12384 23354 12396
rect 25958 12384 25964 12396
rect 26016 12384 26022 12436
rect 22066 12328 22416 12356
rect 18800 12260 19472 12288
rect 18800 12229 18828 12260
rect 19518 12248 19524 12300
rect 19576 12248 19582 12300
rect 20349 12291 20407 12297
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 22186 12288 22192 12300
rect 20395 12260 22192 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 22278 12248 22284 12300
rect 22336 12248 22342 12300
rect 22388 12288 22416 12328
rect 23566 12316 23572 12368
rect 23624 12356 23630 12368
rect 24581 12359 24639 12365
rect 24581 12356 24593 12359
rect 23624 12328 24593 12356
rect 23624 12316 23630 12328
rect 24581 12325 24593 12328
rect 24627 12325 24639 12359
rect 24946 12356 24952 12368
rect 24581 12319 24639 12325
rect 24688 12328 24952 12356
rect 24688 12288 24716 12328
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 22388 12260 24716 12288
rect 24762 12248 24768 12300
rect 24820 12288 24826 12300
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24820 12260 25053 12288
rect 24820 12248 24826 12260
rect 25041 12257 25053 12260
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12257 25191 12291
rect 25133 12251 25191 12257
rect 17788 12192 18736 12220
rect 18785 12223 18843 12229
rect 14384 12124 14780 12152
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 8496 12056 10609 12084
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 10836 12056 10977 12084
rect 10836 12044 10842 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11790 12044 11796 12096
rect 11848 12044 11854 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12342 12084 12348 12096
rect 11940 12056 12348 12084
rect 11940 12044 11946 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 12618 12084 12624 12096
rect 12492 12056 12624 12084
rect 12492 12044 12498 12056
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 12989 12087 13047 12093
rect 12989 12084 13001 12087
rect 12860 12056 13001 12084
rect 12860 12044 12866 12056
rect 12989 12053 13001 12056
rect 13035 12053 13047 12087
rect 12989 12047 13047 12053
rect 13354 12044 13360 12096
rect 13412 12044 13418 12096
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14090 12084 14096 12096
rect 13964 12056 14096 12084
rect 13964 12044 13970 12056
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14366 12044 14372 12096
rect 14424 12044 14430 12096
rect 14752 12084 14780 12124
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 17034 12112 17040 12164
rect 17092 12112 17098 12164
rect 17788 12084 17816 12192
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19536 12220 19564 12248
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19484 12192 19625 12220
rect 19484 12180 19490 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 19518 12112 19524 12164
rect 19576 12152 19582 12164
rect 20088 12152 20116 12183
rect 23658 12180 23664 12232
rect 23716 12180 23722 12232
rect 24946 12180 24952 12232
rect 25004 12180 25010 12232
rect 19576 12124 20116 12152
rect 20732 12124 20838 12152
rect 19576 12112 19582 12124
rect 20732 12096 20760 12124
rect 22554 12112 22560 12164
rect 22612 12112 22618 12164
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 25148 12152 25176 12251
rect 24728 12124 25176 12152
rect 24728 12112 24734 12124
rect 14752 12056 17816 12084
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 17920 12056 18245 12084
rect 17920 12044 17926 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 19337 12087 19395 12093
rect 19337 12053 19349 12087
rect 19383 12084 19395 12087
rect 19429 12087 19487 12093
rect 19429 12084 19441 12087
rect 19383 12056 19441 12084
rect 19383 12053 19395 12056
rect 19337 12047 19395 12053
rect 19429 12053 19441 12056
rect 19475 12084 19487 12087
rect 20714 12084 20720 12096
rect 19475 12056 20720 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 20714 12044 20720 12056
rect 20772 12084 20778 12096
rect 21358 12084 21364 12096
rect 20772 12056 21364 12084
rect 20772 12044 20778 12056
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 21818 12044 21824 12096
rect 21876 12044 21882 12096
rect 23842 12044 23848 12096
rect 23900 12084 23906 12096
rect 24026 12084 24032 12096
rect 23900 12056 24032 12084
rect 23900 12044 23906 12056
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 24394 12044 24400 12096
rect 24452 12084 24458 12096
rect 25593 12087 25651 12093
rect 25593 12084 25605 12087
rect 24452 12056 25605 12084
rect 24452 12044 24458 12056
rect 25593 12053 25605 12056
rect 25639 12053 25651 12087
rect 25593 12047 25651 12053
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2406 11880 2412 11892
rect 2363 11852 2412 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2406 11840 2412 11852
rect 2464 11840 2470 11892
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 2866 11880 2872 11892
rect 2823 11852 2872 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3694 11840 3700 11892
rect 3752 11840 3758 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4801 11883 4859 11889
rect 4801 11880 4813 11883
rect 4764 11852 4813 11880
rect 4764 11840 4770 11852
rect 4801 11849 4813 11852
rect 4847 11849 4859 11883
rect 4801 11843 4859 11849
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5718 11880 5724 11892
rect 5675 11852 5724 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 6052 11852 6745 11880
rect 6052 11840 6058 11852
rect 6733 11849 6745 11852
rect 6779 11849 6791 11883
rect 6733 11843 6791 11849
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8018 11880 8024 11892
rect 7616 11852 8024 11880
rect 7616 11840 7622 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 10502 11840 10508 11892
rect 10560 11840 10566 11892
rect 10965 11883 11023 11889
rect 10965 11849 10977 11883
rect 11011 11880 11023 11883
rect 11882 11880 11888 11892
rect 11011 11852 11888 11880
rect 11011 11849 11023 11852
rect 10965 11843 11023 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 13722 11880 13728 11892
rect 12483 11852 13728 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 13722 11840 13728 11852
rect 13780 11880 13786 11892
rect 16298 11880 16304 11892
rect 13780 11852 16304 11880
rect 13780 11840 13786 11852
rect 16298 11840 16304 11852
rect 16356 11880 16362 11892
rect 16761 11883 16819 11889
rect 16356 11852 16620 11880
rect 16356 11840 16362 11852
rect 7374 11772 7380 11824
rect 7432 11812 7438 11824
rect 7926 11812 7932 11824
rect 7432 11784 7932 11812
rect 7432 11772 7438 11784
rect 7926 11772 7932 11784
rect 7984 11812 7990 11824
rect 7984 11784 8142 11812
rect 7984 11772 7990 11784
rect 9122 11772 9128 11824
rect 9180 11812 9186 11824
rect 9585 11815 9643 11821
rect 9585 11812 9597 11815
rect 9180 11784 9597 11812
rect 9180 11772 9186 11784
rect 9585 11781 9597 11784
rect 9631 11781 9643 11815
rect 10520 11812 10548 11840
rect 11054 11812 11060 11824
rect 10520 11784 11060 11812
rect 9585 11775 9643 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 12345 11815 12403 11821
rect 12345 11812 12357 11815
rect 11624 11784 12357 11812
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2498 11744 2504 11756
rect 1719 11716 2504 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3878 11744 3884 11756
rect 3099 11716 3884 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 5258 11744 5264 11756
rect 4203 11716 5264 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 6546 11744 6552 11756
rect 5767 11716 6552 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5592 11648 5825 11676
rect 5592 11636 5598 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 6086 11676 6092 11688
rect 5859 11648 6092 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6656 11676 6684 11707
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 11624 11753 11652 11784
rect 12345 11781 12357 11784
rect 12391 11781 12403 11815
rect 12345 11775 12403 11781
rect 13446 11772 13452 11824
rect 13504 11772 13510 11824
rect 14458 11772 14464 11824
rect 14516 11772 14522 11824
rect 16592 11812 16620 11852
rect 16761 11849 16773 11883
rect 16807 11880 16819 11883
rect 16850 11880 16856 11892
rect 16807 11852 16856 11880
rect 16807 11849 16819 11852
rect 16761 11843 16819 11849
rect 16850 11840 16856 11852
rect 16908 11880 16914 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 16908 11852 17693 11880
rect 16908 11840 16914 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 35342 11880 35348 11892
rect 17681 11843 17739 11849
rect 18708 11852 35348 11880
rect 16592 11784 16804 11812
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 8996 11716 11621 11744
rect 8996 11704 9002 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 11609 11707 11667 11713
rect 12360 11716 13185 11744
rect 6420 11648 6684 11676
rect 6420 11636 6426 11648
rect 7374 11636 7380 11688
rect 7432 11636 7438 11688
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 8386 11636 8392 11688
rect 8444 11676 8450 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 8444 11648 10333 11676
rect 8444 11636 8450 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 12360 11676 12388 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14792 11716 15393 11744
rect 14792 11704 14798 11716
rect 15381 11713 15393 11716
rect 15427 11744 15439 11747
rect 16666 11744 16672 11756
rect 15427 11716 16672 11744
rect 15427 11713 15439 11716
rect 15381 11707 15439 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16776 11744 16804 11784
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17000 11784 18460 11812
rect 17000 11772 17006 11784
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 16776 11716 17601 11744
rect 17589 11713 17601 11716
rect 17635 11744 17647 11747
rect 17862 11744 17868 11756
rect 17635 11716 17868 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18432 11753 18460 11784
rect 18708 11753 18736 11852
rect 35342 11840 35348 11852
rect 35400 11840 35406 11892
rect 20714 11772 20720 11824
rect 20772 11772 20778 11824
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 21634 11812 21640 11824
rect 21416 11784 21640 11812
rect 21416 11772 21422 11784
rect 21634 11772 21640 11784
rect 21692 11812 21698 11824
rect 21913 11815 21971 11821
rect 21913 11812 21925 11815
rect 21692 11784 21925 11812
rect 21692 11772 21698 11784
rect 21913 11781 21925 11784
rect 21959 11781 21971 11815
rect 21913 11775 21971 11781
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22738 11812 22744 11824
rect 22336 11784 22744 11812
rect 22336 11772 22342 11784
rect 22388 11753 22416 11784
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 23658 11772 23664 11824
rect 23716 11772 23722 11824
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 22373 11747 22431 11753
rect 22373 11713 22385 11747
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 25130 11704 25136 11756
rect 25188 11744 25194 11756
rect 39298 11744 39304 11756
rect 25188 11716 39304 11744
rect 25188 11704 25194 11716
rect 39298 11704 39304 11716
rect 39356 11704 39362 11756
rect 12308 11648 12388 11676
rect 12621 11679 12679 11685
rect 12308 11636 12314 11648
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 3142 11568 3148 11620
rect 3200 11608 3206 11620
rect 7190 11608 7196 11620
rect 3200 11580 7196 11608
rect 3200 11568 3206 11580
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 10686 11608 10692 11620
rect 8720 11580 10692 11608
rect 8720 11568 8726 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 11977 11611 12035 11617
rect 11977 11577 11989 11611
rect 12023 11577 12035 11611
rect 11977 11571 12035 11577
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2866 11540 2872 11552
rect 2004 11512 2872 11540
rect 2004 11500 2010 11512
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3878 11540 3884 11552
rect 3660 11512 3884 11540
rect 3660 11500 3666 11512
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 6638 11540 6644 11552
rect 5307 11512 6644 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 7524 11512 9137 11540
rect 7524 11500 7530 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 11992 11540 12020 11571
rect 12250 11540 12256 11552
rect 11992 11512 12256 11540
rect 9125 11503 9183 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12636 11540 12664 11639
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 16209 11679 16267 11685
rect 13872 11648 14780 11676
rect 13872 11636 13878 11648
rect 14752 11608 14780 11648
rect 16209 11645 16221 11679
rect 16255 11676 16267 11679
rect 16298 11676 16304 11688
rect 16255 11648 16304 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11676 17003 11679
rect 17034 11676 17040 11688
rect 16991 11648 17040 11676
rect 16991 11645 17003 11648
rect 16945 11639 17003 11645
rect 17034 11636 17040 11648
rect 17092 11636 17098 11688
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 17736 11648 17785 11676
rect 17736 11636 17742 11648
rect 17773 11645 17785 11648
rect 17819 11645 17831 11679
rect 17773 11639 17831 11645
rect 19518 11636 19524 11688
rect 19576 11676 19582 11688
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 19576 11648 19717 11676
rect 19576 11636 19582 11648
rect 19705 11645 19717 11648
rect 19751 11645 19763 11679
rect 19705 11639 19763 11645
rect 19978 11636 19984 11688
rect 20036 11636 20042 11688
rect 22649 11679 22707 11685
rect 22649 11645 22661 11679
rect 22695 11676 22707 11679
rect 25866 11676 25872 11688
rect 22695 11648 25872 11676
rect 22695 11645 22707 11648
rect 22649 11639 22707 11645
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 17221 11611 17279 11617
rect 17221 11608 17233 11611
rect 14752 11580 17233 11608
rect 17221 11577 17233 11580
rect 17267 11577 17279 11611
rect 17221 11571 17279 11577
rect 13814 11540 13820 11552
rect 12636 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 13964 11512 14933 11540
rect 13964 11500 13970 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 16390 11540 16396 11552
rect 15252 11512 16396 11540
rect 15252 11500 15258 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 21453 11543 21511 11549
rect 21453 11540 21465 11543
rect 19024 11512 21465 11540
rect 19024 11500 19030 11512
rect 21453 11509 21465 11512
rect 21499 11509 21511 11543
rect 21453 11503 21511 11509
rect 23934 11500 23940 11552
rect 23992 11540 23998 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23992 11512 24133 11540
rect 23992 11500 23998 11512
rect 24121 11509 24133 11512
rect 24167 11509 24179 11543
rect 24121 11503 24179 11509
rect 24394 11500 24400 11552
rect 24452 11540 24458 11552
rect 24581 11543 24639 11549
rect 24581 11540 24593 11543
rect 24452 11512 24593 11540
rect 24452 11500 24458 11512
rect 24581 11509 24593 11512
rect 24627 11509 24639 11543
rect 24581 11503 24639 11509
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3694 11336 3700 11348
rect 2915 11308 3700 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 4028 11308 4169 11336
rect 4028 11296 4034 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 6914 11336 6920 11348
rect 4157 11299 4215 11305
rect 4908 11308 6920 11336
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 3602 11268 3608 11280
rect 3467 11240 3608 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 1854 11160 1860 11212
rect 1912 11160 1918 11212
rect 4908 11144 4936 11308
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7837 11339 7895 11345
rect 7837 11305 7849 11339
rect 7883 11336 7895 11339
rect 8662 11336 8668 11348
rect 7883 11308 8668 11336
rect 7883 11305 7895 11308
rect 7837 11299 7895 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9263 11308 10364 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 7374 11228 7380 11280
rect 7432 11228 7438 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8754 11268 8760 11280
rect 7984 11240 8760 11268
rect 7984 11228 7990 11240
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 9950 11268 9956 11280
rect 9140 11240 9956 11268
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11200 5043 11203
rect 7392 11200 7420 11228
rect 5031 11172 7420 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8076 11172 8401 11200
rect 8076 11160 8082 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 1578 11132 1584 11144
rect 1535 11104 1584 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3237 11135 3295 11141
rect 3237 11132 3249 11135
rect 2832 11104 3249 11132
rect 2832 11092 2838 11104
rect 3237 11101 3249 11104
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4890 11132 4896 11144
rect 4111 11104 4896 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7340 11104 7389 11132
rect 7340 11092 7346 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 9140 11132 9168 11240
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 10336 11268 10364 11308
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13354 11336 13360 11348
rect 12492 11308 13360 11336
rect 12492 11296 12498 11308
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 14182 11296 14188 11348
rect 14240 11296 14246 11348
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 16114 11336 16120 11348
rect 15712 11308 16120 11336
rect 15712 11296 15718 11308
rect 16114 11296 16120 11308
rect 16172 11336 16178 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 16172 11308 16589 11336
rect 16172 11296 16178 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 19242 11336 19248 11348
rect 16577 11299 16635 11305
rect 16684 11308 19248 11336
rect 10336 11240 11744 11268
rect 9306 11160 9312 11212
rect 9364 11200 9370 11212
rect 9769 11203 9827 11209
rect 9769 11200 9781 11203
rect 9364 11172 9781 11200
rect 9364 11160 9370 11172
rect 9769 11169 9781 11172
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11146 11200 11152 11212
rect 11103 11172 11152 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11716 11200 11744 11240
rect 16390 11228 16396 11280
rect 16448 11268 16454 11280
rect 16684 11268 16712 11308
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 23753 11339 23811 11345
rect 23753 11336 23765 11339
rect 20036 11308 23765 11336
rect 20036 11296 20042 11308
rect 23753 11305 23765 11308
rect 23799 11305 23811 11339
rect 23753 11299 23811 11305
rect 16448 11240 16712 11268
rect 16448 11228 16454 11240
rect 18414 11228 18420 11280
rect 18472 11268 18478 11280
rect 18877 11271 18935 11277
rect 18877 11268 18889 11271
rect 18472 11240 18889 11268
rect 18472 11228 18478 11240
rect 18877 11237 18889 11240
rect 18923 11268 18935 11271
rect 18966 11268 18972 11280
rect 18923 11240 18972 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 22646 11228 22652 11280
rect 22704 11228 22710 11280
rect 12250 11200 12256 11212
rect 11716 11172 12256 11200
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13814 11200 13820 11212
rect 13403 11172 13820 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14700 11172 14841 11200
rect 14700 11160 14706 11172
rect 14829 11169 14841 11172
rect 14875 11200 14887 11203
rect 16298 11200 16304 11212
rect 14875 11172 16304 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 17405 11203 17463 11209
rect 16356 11172 17080 11200
rect 16356 11160 16362 11172
rect 17052 11144 17080 11172
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 19242 11200 19248 11212
rect 17451 11172 19248 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 25958 11160 25964 11212
rect 26016 11200 26022 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 26016 11172 29745 11200
rect 26016 11160 26022 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 8343 11104 9168 11132
rect 9585 11135 9643 11141
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 9674 11132 9680 11144
rect 9631 11104 9680 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 10008 11104 10793 11132
rect 10008 11092 10014 11104
rect 10781 11101 10793 11104
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 12952 11104 13921 11132
rect 12952 11092 12958 11104
rect 13909 11101 13921 11104
rect 13955 11132 13967 11135
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 13955 11104 14289 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14277 11101 14289 11104
rect 14323 11132 14335 11135
rect 14366 11132 14372 11144
rect 14323 11104 14372 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14424 11104 14473 11132
rect 14424 11092 14430 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 17092 11104 17141 11132
rect 17092 11092 17098 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11132 20407 11135
rect 20622 11132 20628 11144
rect 20395 11104 20628 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 20622 11092 20628 11104
rect 20680 11132 20686 11144
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 20680 11104 20913 11132
rect 20680 11092 20686 11104
rect 20901 11101 20913 11104
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 23109 11135 23167 11141
rect 23109 11101 23121 11135
rect 23155 11132 23167 11135
rect 24026 11132 24032 11144
rect 23155 11104 24032 11132
rect 23155 11101 23167 11104
rect 23109 11095 23167 11101
rect 24026 11092 24032 11104
rect 24084 11092 24090 11144
rect 31294 11132 31300 11144
rect 31142 11104 31300 11132
rect 31294 11092 31300 11104
rect 31352 11132 31358 11144
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31352 11104 32045 11132
rect 31352 11092 31358 11104
rect 32033 11101 32045 11104
rect 32079 11101 32091 11135
rect 47578 11132 47584 11144
rect 32033 11095 32091 11101
rect 35866 11104 47584 11132
rect 5258 11024 5264 11076
rect 5316 11024 5322 11076
rect 7852 11064 7880 11092
rect 10321 11067 10379 11073
rect 5644 11036 5750 11064
rect 7852 11036 9720 11064
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 4617 10999 4675 11005
rect 4617 10996 4629 10999
rect 3660 10968 4629 10996
rect 3660 10956 3666 10968
rect 4617 10965 4629 10968
rect 4663 10996 4675 10999
rect 5350 10996 5356 11008
rect 4663 10968 5356 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 5350 10956 5356 10968
rect 5408 10996 5414 11008
rect 5644 10996 5672 11036
rect 5408 10968 5672 10996
rect 5408 10956 5414 10968
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 6733 10999 6791 11005
rect 6733 10996 6745 10999
rect 6328 10968 6745 10996
rect 6328 10956 6334 10968
rect 6733 10965 6745 10968
rect 6779 10965 6791 10999
rect 6733 10959 6791 10965
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 9692 11005 9720 11036
rect 10321 11033 10333 11067
rect 10367 11064 10379 11067
rect 10873 11067 10931 11073
rect 10873 11064 10885 11067
rect 10367 11036 10885 11064
rect 10367 11033 10379 11036
rect 10321 11027 10379 11033
rect 10873 11033 10885 11036
rect 10919 11064 10931 11067
rect 11790 11064 11796 11076
rect 10919 11036 11796 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 11882 11024 11888 11076
rect 11940 11024 11946 11076
rect 12618 11024 12624 11076
rect 12676 11024 12682 11076
rect 15105 11067 15163 11073
rect 15105 11033 15117 11067
rect 15151 11064 15163 11067
rect 15194 11064 15200 11076
rect 15151 11036 15200 11064
rect 15151 11033 15163 11036
rect 15105 11027 15163 11033
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 15562 11024 15568 11076
rect 15620 11024 15626 11076
rect 17862 11024 17868 11076
rect 17920 11024 17926 11076
rect 19426 11024 19432 11076
rect 19484 11064 19490 11076
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 19484 11036 19533 11064
rect 19484 11024 19490 11036
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 21634 11024 21640 11076
rect 21692 11024 21698 11076
rect 23658 11024 23664 11076
rect 23716 11064 23722 11076
rect 24121 11067 24179 11073
rect 24121 11064 24133 11067
rect 23716 11036 24133 11064
rect 23716 11024 23722 11036
rect 24121 11033 24133 11036
rect 24167 11064 24179 11067
rect 24394 11064 24400 11076
rect 24167 11036 24400 11064
rect 24167 11033 24179 11036
rect 24121 11027 24179 11033
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 27798 11024 27804 11076
rect 27856 11064 27862 11076
rect 30009 11067 30067 11073
rect 30009 11064 30021 11067
rect 27856 11036 30021 11064
rect 27856 11024 27862 11036
rect 30009 11033 30021 11036
rect 30055 11033 30067 11067
rect 30009 11027 30067 11033
rect 31386 11024 31392 11076
rect 31444 11064 31450 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31444 11036 31769 11064
rect 31444 11024 31450 11036
rect 31757 11033 31769 11036
rect 31803 11064 31815 11067
rect 35866 11064 35894 11104
rect 47578 11092 47584 11104
rect 47636 11092 47642 11144
rect 31803 11036 35894 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 7064 10968 8217 10996
rect 7064 10956 7070 10968
rect 8205 10965 8217 10968
rect 8251 10965 8263 10999
rect 8205 10959 8263 10965
rect 9677 10999 9735 11005
rect 9677 10965 9689 10999
rect 9723 10965 9735 10999
rect 9677 10959 9735 10965
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 13262 10996 13268 11008
rect 9824 10968 13268 10996
rect 9824 10956 9830 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 22094 10956 22100 11008
rect 22152 10996 22158 11008
rect 24302 10996 24308 11008
rect 22152 10968 24308 10996
rect 22152 10956 22158 10968
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1486 10752 1492 10804
rect 1544 10752 1550 10804
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 1854 10792 1860 10804
rect 1811 10764 1860 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 3418 10752 3424 10804
rect 3476 10752 3482 10804
rect 3786 10752 3792 10804
rect 3844 10752 3850 10804
rect 4893 10795 4951 10801
rect 4893 10761 4905 10795
rect 4939 10792 4951 10795
rect 5258 10792 5264 10804
rect 4939 10764 5264 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5960 10764 6009 10792
rect 5960 10752 5966 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6917 10795 6975 10801
rect 6917 10792 6929 10795
rect 6696 10764 6929 10792
rect 6696 10752 6702 10764
rect 6917 10761 6929 10764
rect 6963 10761 6975 10795
rect 6917 10755 6975 10761
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 10137 10795 10195 10801
rect 7248 10764 9352 10792
rect 7248 10752 7254 10764
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2590 10724 2596 10736
rect 2363 10696 2596 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3881 10727 3939 10733
rect 3881 10724 3893 10727
rect 3568 10696 3893 10724
rect 3568 10684 3574 10696
rect 3881 10693 3893 10696
rect 3927 10693 3939 10727
rect 8294 10724 8300 10736
rect 3881 10687 3939 10693
rect 5368 10696 8300 10724
rect 474 10616 480 10668
rect 532 10656 538 10668
rect 934 10656 940 10668
rect 532 10628 940 10656
rect 532 10616 538 10628
rect 934 10616 940 10628
rect 992 10616 998 10668
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 5368 10665 5396 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 8754 10684 8760 10736
rect 8812 10684 8818 10736
rect 9324 10724 9352 10764
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10962 10792 10968 10804
rect 10183 10764 10968 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 11698 10792 11704 10804
rect 11655 10764 11704 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 11793 10795 11851 10801
rect 11793 10761 11805 10795
rect 11839 10792 11851 10795
rect 11974 10792 11980 10804
rect 11839 10764 11980 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12342 10792 12348 10804
rect 12124 10764 12348 10792
rect 12124 10752 12130 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13170 10792 13176 10804
rect 12728 10764 13176 10792
rect 12728 10736 12756 10764
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 13262 10752 13268 10804
rect 13320 10792 13326 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 13320 10764 14381 10792
rect 13320 10752 13326 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 14826 10752 14832 10804
rect 14884 10752 14890 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 15804 10764 16865 10792
rect 15804 10752 15810 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 19518 10792 19524 10804
rect 16853 10755 16911 10761
rect 17512 10764 19524 10792
rect 10781 10727 10839 10733
rect 10781 10724 10793 10727
rect 9324 10696 10793 10724
rect 10781 10693 10793 10696
rect 10827 10693 10839 10727
rect 10781 10687 10839 10693
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 12710 10724 12716 10736
rect 10928 10696 12716 10724
rect 10928 10684 10934 10696
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 12894 10684 12900 10736
rect 12952 10684 12958 10736
rect 14458 10684 14464 10736
rect 14516 10724 14522 10736
rect 15933 10727 15991 10733
rect 15933 10724 15945 10727
rect 14516 10696 15945 10724
rect 14516 10684 14522 10696
rect 15933 10693 15945 10696
rect 15979 10693 15991 10727
rect 15933 10687 15991 10693
rect 16025 10727 16083 10733
rect 16025 10693 16037 10727
rect 16071 10724 16083 10727
rect 17218 10724 17224 10736
rect 16071 10696 17224 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 2133 10659 2191 10665
rect 2133 10656 2145 10659
rect 1912 10628 2145 10656
rect 1912 10616 1918 10628
rect 2133 10625 2145 10628
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 2792 10452 2820 10619
rect 4264 10588 4292 10619
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6328 10628 7144 10656
rect 6328 10616 6334 10628
rect 5442 10588 5448 10600
rect 4264 10560 5448 10588
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 7116 10597 7144 10628
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9640 10628 11008 10656
rect 9640 10616 9646 10628
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 7024 10520 7052 10551
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7432 10560 7757 10588
rect 7432 10548 7438 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8021 10591 8079 10597
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8570 10588 8576 10600
rect 8067 10560 8576 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 5132 10492 7052 10520
rect 5132 10480 5138 10492
rect 6270 10452 6276 10464
rect 2792 10424 6276 10452
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6638 10452 6644 10464
rect 6595 10424 6644 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 7760 10452 7788 10551
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 9030 10548 9036 10600
rect 9088 10588 9094 10600
rect 10980 10597 11008 10628
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 11664 10628 12173 10656
rect 11664 10616 11670 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 16942 10656 16948 10668
rect 14844 10628 16948 10656
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9088 10560 9781 10588
rect 9088 10548 9094 10560
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 10873 10591 10931 10597
rect 10873 10557 10885 10591
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10557 11023 10591
rect 10965 10551 11023 10557
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 13722 10588 13728 10600
rect 12483 10560 13728 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 10042 10520 10048 10532
rect 9180 10492 10048 10520
rect 9180 10480 9186 10492
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 10888 10520 10916 10551
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 11974 10520 11980 10532
rect 10888 10492 11980 10520
rect 11974 10480 11980 10492
rect 12032 10480 12038 10532
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 14844 10520 14872 10628
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17512 10665 17540 10764
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 21453 10795 21511 10801
rect 21453 10792 21465 10795
rect 19628 10764 21465 10792
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 19628 10724 19656 10764
rect 21453 10761 21465 10764
rect 21499 10761 21511 10795
rect 21453 10755 21511 10761
rect 21634 10752 21640 10804
rect 21692 10792 21698 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 21692 10764 21833 10792
rect 21692 10752 21698 10764
rect 21821 10761 21833 10764
rect 21867 10761 21879 10795
rect 21821 10755 21879 10761
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 22612 10764 22845 10792
rect 22612 10752 22618 10764
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 22833 10755 22891 10761
rect 21266 10724 21272 10736
rect 17920 10696 18262 10724
rect 19168 10696 19656 10724
rect 21206 10696 21272 10724
rect 17920 10684 17926 10696
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17184 10628 17509 10656
rect 17184 10616 17190 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 16114 10588 16120 10600
rect 15059 10560 16120 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 13596 10492 14872 10520
rect 15565 10523 15623 10529
rect 13596 10480 13602 10492
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 15930 10520 15936 10532
rect 15611 10492 15936 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 8386 10452 8392 10464
rect 7760 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 10410 10412 10416 10464
rect 10468 10412 10474 10464
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 12618 10452 12624 10464
rect 12216 10424 12624 10452
rect 12216 10412 12222 10424
rect 12618 10412 12624 10424
rect 12676 10452 12682 10464
rect 12894 10452 12900 10464
rect 12676 10424 12900 10452
rect 12676 10412 12682 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13228 10424 13921 10452
rect 13228 10412 13234 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 16224 10452 16252 10551
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 16356 10560 17785 10588
rect 16356 10548 16362 10560
rect 17773 10557 17785 10560
rect 17819 10588 17831 10591
rect 19058 10588 19064 10600
rect 17819 10560 19064 10588
rect 17819 10557 17831 10560
rect 17773 10551 17831 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 18874 10480 18880 10532
rect 18932 10520 18938 10532
rect 19168 10520 19196 10696
rect 21266 10684 21272 10696
rect 21324 10724 21330 10736
rect 21652 10724 21680 10752
rect 21324 10696 21680 10724
rect 21324 10684 21330 10696
rect 21818 10616 21824 10668
rect 21876 10656 21882 10668
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21876 10628 22201 10656
rect 21876 10616 21882 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 22704 10628 23305 10656
rect 22704 10616 22710 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 19981 10591 20039 10597
rect 19751 10560 19840 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 18932 10492 19196 10520
rect 18932 10480 18938 10492
rect 18414 10452 18420 10464
rect 16224 10424 18420 10452
rect 13909 10415 13967 10421
rect 18414 10412 18420 10424
rect 18472 10452 18478 10464
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 18472 10424 19257 10452
rect 18472 10412 18478 10424
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 19812 10452 19840 10560
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 20027 10560 23949 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 20622 10452 20628 10464
rect 19576 10424 20628 10452
rect 19576 10412 19582 10424
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 24302 10412 24308 10464
rect 24360 10452 24366 10464
rect 34882 10452 34888 10464
rect 24360 10424 34888 10452
rect 24360 10412 24366 10424
rect 34882 10412 34888 10424
rect 34940 10412 34946 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 382 10208 388 10260
rect 440 10248 446 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 440 10220 3065 10248
rect 440 10208 446 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 3602 10208 3608 10260
rect 3660 10208 3666 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4120 10220 4169 10248
rect 4120 10208 4126 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 4580 10220 6193 10248
rect 4580 10208 4586 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6641 10251 6699 10257
rect 6641 10248 6653 10251
rect 6604 10220 6653 10248
rect 6604 10208 6610 10220
rect 6641 10217 6653 10220
rect 6687 10217 6699 10251
rect 13538 10248 13544 10260
rect 6641 10211 6699 10217
rect 6748 10220 13544 10248
rect 6748 10180 6776 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13630 10208 13636 10260
rect 13688 10208 13694 10260
rect 16666 10208 16672 10260
rect 16724 10208 16730 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 17276 10220 18889 10248
rect 17276 10208 17282 10220
rect 18877 10217 18889 10220
rect 18923 10248 18935 10251
rect 20162 10248 20168 10260
rect 18923 10220 20168 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22244 10220 22385 10248
rect 22244 10208 22250 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 22373 10211 22431 10217
rect 5920 10152 6776 10180
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1452 10084 1593 10112
rect 1452 10072 1458 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1026 10004 1032 10056
rect 1084 10044 1090 10056
rect 1857 10047 1915 10053
rect 1857 10044 1869 10047
rect 1084 10016 1869 10044
rect 1084 10004 1090 10016
rect 1857 10013 1869 10016
rect 1903 10013 1915 10047
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 1857 10007 1915 10013
rect 2746 10016 4997 10044
rect 290 9868 296 9920
rect 348 9908 354 9920
rect 2746 9908 2774 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 2958 9936 2964 9988
rect 3016 9936 3022 9988
rect 4062 9936 4068 9988
rect 4120 9936 4126 9988
rect 4801 9979 4859 9985
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 5258 9976 5264 9988
rect 4847 9948 5264 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5258 9936 5264 9948
rect 5316 9976 5322 9988
rect 5920 9976 5948 10152
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 13909 10183 13967 10189
rect 7524 10152 8432 10180
rect 7524 10140 7530 10152
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 6052 10084 7205 10112
rect 6052 10072 6058 10084
rect 7193 10081 7205 10084
rect 7239 10081 7251 10115
rect 7193 10075 7251 10081
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 8404 10121 8432 10152
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 14366 10180 14372 10192
rect 13955 10152 14372 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 16390 10140 16396 10192
rect 16448 10140 16454 10192
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 7800 10084 8309 10112
rect 7800 10072 7806 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 9858 10112 9864 10124
rect 8389 10075 8447 10081
rect 8496 10084 9864 10112
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 8496 10044 8524 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 14642 10112 14648 10124
rect 11440 10084 14648 10112
rect 11440 10053 11468 10084
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 16298 10112 16304 10124
rect 14976 10084 16304 10112
rect 14976 10072 14982 10084
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17126 10112 17132 10124
rect 16908 10084 17132 10112
rect 16908 10072 16914 10084
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 19518 10072 19524 10124
rect 19576 10072 19582 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10112 19855 10115
rect 22646 10112 22652 10124
rect 19843 10084 22652 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 22646 10072 22652 10084
rect 22704 10072 22710 10124
rect 7147 10016 8524 10044
rect 9125 10047 9183 10053
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 21266 10044 21272 10056
rect 20930 10016 21272 10044
rect 11425 10007 11483 10013
rect 5316 9948 5948 9976
rect 5316 9936 5322 9948
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9140 9976 9168 10007
rect 8444 9948 9168 9976
rect 8444 9936 8450 9948
rect 9398 9936 9404 9988
rect 9456 9936 9462 9988
rect 9858 9936 9864 9988
rect 9916 9936 9922 9988
rect 11440 9976 11468 10007
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 21726 10004 21732 10056
rect 21784 10044 21790 10056
rect 24670 10044 24676 10056
rect 21784 10016 24676 10044
rect 21784 10004 21790 10016
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 11606 9976 11612 9988
rect 11440 9948 11612 9976
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9976 11759 9979
rect 11790 9976 11796 9988
rect 11747 9948 11796 9976
rect 11747 9945 11759 9948
rect 11701 9939 11759 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 12158 9976 12164 9988
rect 12084 9948 12164 9976
rect 348 9880 2774 9908
rect 348 9868 354 9880
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7009 9911 7067 9917
rect 7009 9908 7021 9911
rect 6972 9880 7021 9908
rect 6972 9868 6978 9880
rect 7009 9877 7021 9880
rect 7055 9877 7067 9911
rect 7009 9871 7067 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7800 9880 7849 9908
rect 7800 9868 7806 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 10318 9908 10324 9920
rect 8251 9880 10324 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 10870 9868 10876 9920
rect 10928 9868 10934 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11974 9908 11980 9920
rect 11204 9880 11980 9908
rect 11204 9868 11210 9880
rect 11974 9868 11980 9880
rect 12032 9908 12038 9920
rect 12084 9908 12112 9948
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 14921 9979 14979 9985
rect 14921 9945 14933 9979
rect 14967 9976 14979 9979
rect 15194 9976 15200 9988
rect 14967 9948 15200 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15304 9948 15410 9976
rect 12032 9880 12112 9908
rect 12032 9868 12038 9880
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 12768 9880 13185 9908
rect 12768 9868 12774 9880
rect 13173 9877 13185 9880
rect 13219 9877 13231 9911
rect 13173 9871 13231 9877
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13320 9880 13461 9908
rect 13320 9868 13326 9880
rect 13449 9877 13461 9880
rect 13495 9908 13507 9911
rect 13630 9908 13636 9920
rect 13495 9880 13636 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13630 9868 13636 9880
rect 13688 9908 13694 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13688 9880 14105 9908
rect 13688 9868 13694 9880
rect 14093 9877 14105 9880
rect 14139 9908 14151 9911
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 14139 9880 14289 9908
rect 14139 9877 14151 9880
rect 14093 9871 14151 9877
rect 14277 9877 14289 9880
rect 14323 9908 14335 9911
rect 15304 9908 15332 9948
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 17862 9976 17868 9988
rect 17788 9948 17868 9976
rect 15562 9908 15568 9920
rect 14323 9880 15568 9908
rect 14323 9877 14335 9880
rect 14277 9871 14335 9877
rect 15562 9868 15568 9880
rect 15620 9908 15626 9920
rect 17788 9908 17816 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 18690 9908 18696 9920
rect 15620 9880 18696 9908
rect 15620 9868 15626 9880
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 9306 9704 9312 9716
rect 3252 9676 3464 9704
rect 1486 9596 1492 9648
rect 1544 9596 1550 9648
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1765 9639 1823 9645
rect 1765 9636 1777 9639
rect 1728 9608 1777 9636
rect 1728 9596 1734 9608
rect 1765 9605 1777 9608
rect 1811 9605 1823 9639
rect 1765 9599 1823 9605
rect 2130 9596 2136 9648
rect 2188 9596 2194 9648
rect 2148 9568 2176 9596
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2148 9540 2421 9568
rect 2409 9537 2421 9540
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 3252 9500 3280 9676
rect 3326 9596 3332 9648
rect 3384 9596 3390 9648
rect 3436 9636 3464 9676
rect 7852 9676 9312 9704
rect 4246 9636 4252 9648
rect 3436 9608 4252 9636
rect 4246 9596 4252 9608
rect 4304 9636 4310 9648
rect 5074 9636 5080 9648
rect 4304 9608 5080 9636
rect 4304 9596 4310 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5994 9596 6000 9648
rect 6052 9596 6058 9648
rect 7006 9636 7012 9648
rect 6104 9608 7012 9636
rect 3418 9568 3424 9580
rect 2179 9472 3280 9500
rect 3344 9540 3424 9568
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 3344 9432 3372 9540
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3936 9540 4077 9568
rect 3936 9528 3942 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4172 9540 5120 9568
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 4172 9500 4200 9540
rect 3743 9472 4200 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 4246 9460 4252 9512
rect 4304 9460 4310 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 5092 9500 5120 9540
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5224 9540 5365 9568
rect 5224 9528 5230 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 6104 9568 6132 9608
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 7285 9571 7343 9577
rect 5500 9540 6132 9568
rect 6564 9540 7236 9568
rect 5500 9528 5506 9540
rect 6564 9500 6592 9540
rect 5092 9472 6592 9500
rect 6641 9503 6699 9509
rect 4709 9463 4767 9469
rect 6641 9469 6653 9503
rect 6687 9469 6699 9503
rect 7208 9500 7236 9540
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7852 9568 7880 9676
rect 9306 9664 9312 9676
rect 9364 9704 9370 9716
rect 10502 9704 10508 9716
rect 9364 9676 10508 9704
rect 9364 9664 9370 9676
rect 10502 9664 10508 9676
rect 10560 9704 10566 9716
rect 10870 9704 10876 9716
rect 10560 9676 10876 9704
rect 10560 9664 10566 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11146 9704 11152 9716
rect 10980 9676 11152 9704
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8665 9639 8723 9645
rect 8665 9636 8677 9639
rect 7975 9608 8677 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8665 9605 8677 9608
rect 8711 9605 8723 9639
rect 8665 9599 8723 9605
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 8938 9636 8944 9648
rect 8812 9608 8944 9636
rect 8812 9596 8818 9608
rect 8938 9596 8944 9608
rect 8996 9636 9002 9648
rect 8996 9608 9154 9636
rect 8996 9596 9002 9608
rect 10686 9596 10692 9648
rect 10744 9596 10750 9648
rect 10980 9636 11008 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 14274 9704 14280 9716
rect 11716 9676 14280 9704
rect 11716 9636 11744 9676
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 21545 9707 21603 9713
rect 21545 9704 21557 9707
rect 21416 9676 21557 9704
rect 21416 9664 21422 9676
rect 21545 9673 21557 9676
rect 21591 9673 21603 9707
rect 21545 9667 21603 9673
rect 22738 9664 22744 9716
rect 22796 9704 22802 9716
rect 24578 9704 24584 9716
rect 22796 9676 24584 9704
rect 22796 9664 22802 9676
rect 24578 9664 24584 9676
rect 24636 9664 24642 9716
rect 10888 9608 11008 9636
rect 11072 9608 11744 9636
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 7331 9540 7880 9568
rect 9876 9540 10425 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 9876 9512 9904 9540
rect 10413 9537 10425 9540
rect 10459 9568 10471 9571
rect 10888 9568 10916 9608
rect 10459 9540 10916 9568
rect 10965 9571 11023 9577
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11072 9568 11100 9608
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12032 9608 12466 9636
rect 12032 9596 12038 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13725 9639 13783 9645
rect 13725 9636 13737 9639
rect 13688 9608 13737 9636
rect 13688 9596 13694 9608
rect 13725 9605 13737 9608
rect 13771 9605 13783 9639
rect 15102 9636 15108 9648
rect 13725 9599 13783 9605
rect 13832 9608 15108 9636
rect 11011 9540 11100 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11664 9540 11713 9568
rect 11664 9528 11670 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 13832 9568 13860 9608
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 15562 9596 15568 9648
rect 15620 9596 15626 9648
rect 17129 9639 17187 9645
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 17218 9636 17224 9648
rect 17175 9608 17224 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 18690 9636 18696 9648
rect 18354 9608 18696 9636
rect 18690 9596 18696 9608
rect 18748 9596 18754 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 19567 9608 20852 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 13320 9540 13860 9568
rect 13320 9528 13326 9540
rect 14550 9528 14556 9580
rect 14608 9528 14614 9580
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 18564 9540 19441 9568
rect 18564 9528 18570 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19429 9531 19487 9537
rect 19536 9540 20269 9568
rect 8294 9500 8300 9512
rect 7208 9472 8300 9500
rect 6641 9463 6699 9469
rect 2648 9404 3372 9432
rect 2648 9392 2654 9404
rect 3418 9392 3424 9444
rect 3476 9392 3482 9444
rect 1670 9324 1676 9376
rect 1728 9324 1734 9376
rect 3878 9324 3884 9376
rect 3936 9324 3942 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4724 9364 4752 9463
rect 6656 9432 6684 9463
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8386 9460 8392 9512
rect 8444 9460 8450 9512
rect 8496 9472 9720 9500
rect 8496 9432 8524 9472
rect 6656 9404 8524 9432
rect 6914 9364 6920 9376
rect 4663 9336 6920 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 9692 9364 9720 9472
rect 9858 9460 9864 9512
rect 9916 9460 9922 9512
rect 11146 9500 11152 9512
rect 9968 9472 11152 9500
rect 9968 9364 9996 9472
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11974 9460 11980 9512
rect 12032 9460 12038 9512
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 12400 9472 13461 9500
rect 12400 9460 12406 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14182 9500 14188 9512
rect 14047 9472 14188 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 14826 9460 14832 9512
rect 14884 9460 14890 9512
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15436 9472 16313 9500
rect 15436 9460 15442 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16408 9472 18736 9500
rect 11698 9432 11704 9444
rect 10152 9404 11704 9432
rect 9692 9336 9996 9364
rect 10042 9324 10048 9376
rect 10100 9364 10106 9376
rect 10152 9373 10180 9404
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 14108 9404 14320 9432
rect 10137 9367 10195 9373
rect 10137 9364 10149 9367
rect 10100 9336 10149 9364
rect 10100 9324 10106 9336
rect 10137 9333 10149 9336
rect 10183 9333 10195 9367
rect 10137 9327 10195 9333
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 14108 9364 14136 9404
rect 10928 9336 14136 9364
rect 10928 9324 10934 9336
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 14292 9364 14320 9404
rect 16408 9364 16436 9472
rect 14292 9336 16436 9364
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 17368 9336 18613 9364
rect 17368 9324 17374 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18708 9364 18736 9472
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19536 9500 19564 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20824 9568 20852 9608
rect 20898 9596 20904 9648
rect 20956 9596 20962 9648
rect 22094 9636 22100 9648
rect 21008 9608 22100 9636
rect 21008 9568 21036 9608
rect 22094 9596 22100 9608
rect 22152 9596 22158 9648
rect 22646 9596 22652 9648
rect 22704 9596 22710 9648
rect 27798 9596 27804 9648
rect 27856 9596 27862 9648
rect 20824 9540 21036 9568
rect 20257 9531 20315 9537
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 23934 9568 23940 9580
rect 22060 9540 23940 9568
rect 22060 9528 22066 9540
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 24084 9540 27169 9568
rect 24084 9528 24090 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 19024 9472 19564 9500
rect 19705 9503 19763 9509
rect 19024 9460 19030 9472
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 21266 9500 21272 9512
rect 19751 9472 21272 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 19061 9435 19119 9441
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 26050 9432 26056 9444
rect 19107 9404 26056 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 26050 9392 26056 9404
rect 26108 9392 26114 9444
rect 19150 9364 19156 9376
rect 18708 9336 19156 9364
rect 18601 9327 18659 9333
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1452 9132 1593 9160
rect 1452 9120 1458 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2038 9120 2044 9172
rect 2096 9120 2102 9172
rect 4706 9120 4712 9172
rect 4764 9120 4770 9172
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4948 9132 4997 9160
rect 4948 9120 4954 9132
rect 4985 9129 4997 9132
rect 5031 9129 5043 9163
rect 6178 9160 6184 9172
rect 4985 9123 5043 9129
rect 5460 9132 6184 9160
rect 1670 9052 1676 9104
rect 1728 9092 1734 9104
rect 2498 9092 2504 9104
rect 1728 9064 2504 9092
rect 1728 9052 1734 9064
rect 2498 9052 2504 9064
rect 2556 9092 2562 9104
rect 5460 9092 5488 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6270 9120 6276 9172
rect 6328 9120 6334 9172
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7650 9160 7656 9172
rect 7423 9132 7656 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10192 9132 10425 9160
rect 10192 9120 10198 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 13354 9160 13360 9172
rect 10413 9123 10471 9129
rect 11624 9132 13360 9160
rect 7466 9092 7472 9104
rect 2556 9064 5488 9092
rect 5552 9064 7472 9092
rect 2556 9052 2562 9064
rect 1210 8984 1216 9036
rect 1268 9024 1274 9036
rect 2593 9027 2651 9033
rect 1268 8996 1900 9024
rect 1268 8984 1274 8996
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 1872 8956 1900 8996
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 5552 9024 5580 9064
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 8754 9092 8760 9104
rect 8496 9064 8760 9092
rect 7098 9024 7104 9036
rect 2639 8996 5580 9024
rect 5644 8996 7104 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 1872 8928 2881 8956
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 4028 8928 4077 8956
rect 4028 8916 4034 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5350 8956 5356 8968
rect 5224 8928 5356 8956
rect 5224 8916 5230 8928
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5644 8965 5672 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8496 9033 8524 9064
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 9582 9092 9588 9104
rect 8812 9064 9588 9092
rect 8812 9052 8818 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 9953 9095 10011 9101
rect 9953 9061 9965 9095
rect 9999 9092 10011 9095
rect 11624 9092 11652 9132
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 15028 9132 17724 9160
rect 9999 9064 11652 9092
rect 14369 9095 14427 9101
rect 9999 9061 10011 9064
rect 9953 9055 10011 9061
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 14415 9064 14964 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 7892 8996 8309 9024
rect 7892 8984 7898 8996
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 10318 9024 10324 9036
rect 8481 8987 8539 8993
rect 9324 8996 10324 9024
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7708 8928 8217 8956
rect 7708 8916 7714 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 8938 8956 8944 8968
rect 8720 8928 8944 8956
rect 8720 8916 8726 8928
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9324 8965 9352 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10686 8956 10692 8968
rect 10192 8928 10692 8956
rect 10192 8916 10198 8928
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10870 8916 10876 8968
rect 10928 8916 10934 8968
rect 10980 8956 11008 8987
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 11756 8996 12173 9024
rect 11756 8984 11762 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 12897 9027 12955 9033
rect 12897 9024 12909 9027
rect 12860 8996 12909 9024
rect 12860 8984 12866 8996
rect 12897 8993 12909 8996
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13906 9024 13912 9036
rect 13412 8996 13912 9024
rect 13412 8984 13418 8996
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 12710 8956 12716 8968
rect 10980 8928 12716 8956
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 4246 8848 4252 8900
rect 4304 8848 4310 8900
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 8478 8888 8484 8900
rect 4396 8860 8484 8888
rect 4396 8848 4402 8860
rect 8478 8848 8484 8860
rect 8536 8848 8542 8900
rect 9582 8888 9588 8900
rect 8956 8860 9588 8888
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2498 8820 2504 8832
rect 2363 8792 2504 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2498 8780 2504 8792
rect 2556 8820 2562 8832
rect 2682 8820 2688 8832
rect 2556 8792 2688 8820
rect 2556 8780 2562 8792
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 7374 8820 7380 8832
rect 5224 8792 7380 8820
rect 5224 8780 5230 8792
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 8956 8820 8984 8860
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 9916 8860 11989 8888
rect 9916 8848 9922 8860
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 12069 8891 12127 8897
rect 12069 8857 12081 8891
rect 12115 8888 12127 8891
rect 12158 8888 12164 8900
rect 12115 8860 12164 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 14182 8888 14188 8900
rect 12308 8860 14188 8888
rect 12308 8848 12314 8860
rect 14182 8848 14188 8860
rect 14240 8888 14246 8900
rect 14829 8891 14887 8897
rect 14829 8888 14841 8891
rect 14240 8860 14841 8888
rect 14240 8848 14246 8860
rect 14829 8857 14841 8860
rect 14875 8857 14887 8891
rect 14936 8888 14964 9064
rect 15028 9033 15056 9132
rect 15562 9052 15568 9104
rect 15620 9092 15626 9104
rect 15657 9095 15715 9101
rect 15657 9092 15669 9095
rect 15620 9064 15669 9092
rect 15620 9052 15626 9064
rect 15657 9061 15669 9064
rect 15703 9061 15715 9095
rect 17696 9092 17724 9132
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 18877 9163 18935 9169
rect 18877 9160 18889 9163
rect 17828 9132 18889 9160
rect 17828 9120 17834 9132
rect 18877 9129 18889 9132
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 19426 9120 19432 9172
rect 19484 9120 19490 9172
rect 20993 9163 21051 9169
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 21174 9160 21180 9172
rect 21039 9132 21180 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 27893 9163 27951 9169
rect 27893 9129 27905 9163
rect 27939 9160 27951 9163
rect 28721 9163 28779 9169
rect 28721 9160 28733 9163
rect 27939 9132 28733 9160
rect 27939 9129 27951 9132
rect 27893 9123 27951 9129
rect 28721 9129 28733 9132
rect 28767 9160 28779 9163
rect 31386 9160 31392 9172
rect 28767 9132 31392 9160
rect 28767 9129 28779 9132
rect 28721 9123 28779 9129
rect 31386 9120 31392 9132
rect 31444 9120 31450 9172
rect 21726 9092 21732 9104
rect 17696 9064 21732 9092
rect 15657 9055 15715 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 15013 9027 15071 9033
rect 15013 8993 15025 9027
rect 15059 8993 15071 9027
rect 15013 8987 15071 8993
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16850 9024 16856 9036
rect 16071 8996 16856 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 24762 8984 24768 9036
rect 24820 9024 24826 9036
rect 35434 9024 35440 9036
rect 24820 8996 35440 9024
rect 24820 8984 24826 8996
rect 35434 8984 35440 8996
rect 35492 8984 35498 9036
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 21266 8956 21272 8968
rect 20395 8928 21272 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8956 27675 8959
rect 27663 8928 28580 8956
rect 27663 8925 27675 8928
rect 27617 8919 27675 8925
rect 16301 8891 16359 8897
rect 14936 8860 16252 8888
rect 14829 8851 14887 8857
rect 7883 8792 8984 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 9088 8792 10793 8820
rect 9088 8780 9094 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 10781 8783 10839 8789
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11330 8820 11336 8832
rect 10928 8792 11336 8820
rect 10928 8780 10934 8792
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 11790 8820 11796 8832
rect 11655 8792 11796 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13630 8820 13636 8832
rect 12584 8792 13636 8820
rect 12584 8780 12590 8792
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 15102 8820 15108 8832
rect 14783 8792 15108 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16224 8820 16252 8860
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 16574 8888 16580 8900
rect 16347 8860 16580 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 16758 8848 16764 8900
rect 16816 8848 16822 8900
rect 20530 8888 20536 8900
rect 17604 8860 20536 8888
rect 17604 8820 17632 8860
rect 20530 8848 20536 8860
rect 20588 8848 20594 8900
rect 16224 8792 17632 8820
rect 17770 8780 17776 8832
rect 17828 8780 17834 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19705 8823 19763 8829
rect 19705 8820 19717 8823
rect 19576 8792 19717 8820
rect 19576 8780 19582 8792
rect 19705 8789 19717 8792
rect 19751 8820 19763 8823
rect 19889 8823 19947 8829
rect 19889 8820 19901 8823
rect 19751 8792 19901 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19889 8789 19901 8792
rect 19935 8789 19947 8823
rect 19889 8783 19947 8789
rect 26234 8780 26240 8832
rect 26292 8820 26298 8832
rect 28552 8829 28580 8928
rect 28077 8823 28135 8829
rect 28077 8820 28089 8823
rect 26292 8792 28089 8820
rect 26292 8780 26298 8792
rect 28077 8789 28089 8792
rect 28123 8789 28135 8823
rect 28077 8783 28135 8789
rect 28537 8823 28595 8829
rect 28537 8789 28549 8823
rect 28583 8820 28595 8823
rect 28718 8820 28724 8832
rect 28583 8792 28724 8820
rect 28583 8789 28595 8792
rect 28537 8783 28595 8789
rect 28718 8780 28724 8792
rect 28776 8780 28782 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1762 8616 1768 8628
rect 1627 8588 1768 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 4798 8616 4804 8628
rect 1964 8588 4804 8616
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 1854 8480 1860 8492
rect 1811 8452 1860 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 1964 8412 1992 8588
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5767 8588 5825 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5813 8585 5825 8588
rect 5859 8616 5871 8619
rect 5902 8616 5908 8628
rect 5859 8588 5908 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 9674 8616 9680 8628
rect 6236 8588 9680 8616
rect 6236 8576 6242 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9858 8576 9864 8628
rect 9916 8576 9922 8628
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10410 8616 10416 8628
rect 10275 8588 10416 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11054 8576 11060 8628
rect 11112 8576 11118 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11606 8576 11612 8628
rect 11664 8576 11670 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12802 8616 12808 8628
rect 11931 8588 12808 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 14366 8576 14372 8628
rect 14424 8576 14430 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16482 8616 16488 8628
rect 16347 8588 16488 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16574 8576 16580 8628
rect 16632 8616 16638 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 16632 8588 17877 8616
rect 16632 8576 16638 8588
rect 17865 8585 17877 8588
rect 17911 8585 17923 8619
rect 17865 8579 17923 8585
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18690 8616 18696 8628
rect 18279 8588 18696 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19242 8576 19248 8628
rect 19300 8576 19306 8628
rect 2038 8508 2044 8560
rect 2096 8548 2102 8560
rect 4338 8548 4344 8560
rect 2096 8520 2452 8548
rect 2096 8508 2102 8520
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 2424 8480 2452 8520
rect 2746 8520 4344 8548
rect 2746 8480 2774 8520
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 5994 8548 6000 8560
rect 4672 8520 6000 8548
rect 4672 8508 4678 8520
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 6270 8508 6276 8560
rect 6328 8548 6334 8560
rect 6328 8520 8294 8548
rect 6328 8508 6334 8520
rect 2424 8452 2774 8480
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 3476 8452 3617 8480
rect 3476 8440 3482 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 6549 8483 6607 8489
rect 5040 8452 5580 8480
rect 5040 8440 5046 8452
rect 2041 8415 2099 8421
rect 2041 8412 2053 8415
rect 1964 8384 2053 8412
rect 2041 8381 2053 8384
rect 2087 8381 2099 8415
rect 2041 8375 2099 8381
rect 2130 8372 2136 8424
rect 2188 8412 2194 8424
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 2188 8384 3341 8412
rect 2188 8372 2194 8384
rect 3329 8381 3341 8384
rect 3375 8381 3387 8415
rect 3329 8375 3387 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4571 8384 4629 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 4617 8381 4629 8384
rect 4663 8412 4675 8415
rect 5442 8412 5448 8424
rect 4663 8384 5448 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 5552 8412 5580 8452
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6730 8480 6736 8492
rect 6595 8452 6736 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7616 8452 7941 8480
rect 7616 8440 7622 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 8266 8480 8294 8520
rect 9398 8508 9404 8560
rect 9456 8508 9462 8560
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 10321 8551 10379 8557
rect 10321 8548 10333 8551
rect 9640 8520 10333 8548
rect 9640 8508 9646 8520
rect 10321 8517 10333 8520
rect 10367 8517 10379 8551
rect 10321 8511 10379 8517
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 10560 8520 10640 8548
rect 10560 8508 10566 8520
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8266 8452 8493 8480
rect 7929 8443 7987 8449
rect 8481 8449 8493 8452
rect 8527 8480 8539 8483
rect 8662 8480 8668 8492
rect 8527 8452 8668 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 5552 8384 6837 8412
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 7834 8412 7840 8424
rect 7708 8384 7840 8412
rect 7708 8372 7714 8384
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8110 8372 8116 8424
rect 8168 8372 8174 8424
rect 9858 8412 9864 8424
rect 8220 8384 9864 8412
rect 3142 8304 3148 8356
rect 3200 8344 3206 8356
rect 6638 8344 6644 8356
rect 3200 8316 6644 8344
rect 3200 8304 3206 8316
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 8220 8344 8248 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10505 8415 10563 8421
rect 10505 8381 10517 8415
rect 10551 8412 10563 8415
rect 10612 8412 10640 8520
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 12253 8551 12311 8557
rect 12253 8548 12265 8551
rect 11480 8520 12265 8548
rect 11480 8508 11486 8520
rect 12253 8517 12265 8520
rect 12299 8517 12311 8551
rect 12253 8511 12311 8517
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 12584 8520 14841 8548
rect 12584 8508 12590 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 22002 8548 22008 8560
rect 14829 8511 14887 8517
rect 15580 8520 22008 8548
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 12084 8452 12357 8480
rect 12084 8412 12112 8452
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 14182 8480 14188 8492
rect 13495 8452 14188 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14332 8452 14749 8480
rect 14332 8440 14338 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 15580 8480 15608 8520
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 14737 8443 14795 8449
rect 14844 8452 15608 8480
rect 10551 8384 10640 8412
rect 10796 8384 12112 8412
rect 12529 8415 12587 8421
rect 10551 8381 10563 8384
rect 10505 8375 10563 8381
rect 7616 8316 8248 8344
rect 7616 8304 7622 8316
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 10796 8344 10824 8384
rect 12529 8381 12541 8415
rect 12575 8412 12587 8415
rect 12575 8384 13032 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 8352 8316 10824 8344
rect 10965 8347 11023 8353
rect 8352 8304 8358 8316
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11054 8344 11060 8356
rect 11011 8316 11060 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11606 8304 11612 8356
rect 11664 8344 11670 8356
rect 12342 8344 12348 8356
rect 11664 8316 12348 8344
rect 11664 8304 11670 8316
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 5353 8279 5411 8285
rect 5353 8245 5365 8279
rect 5399 8276 5411 8279
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5399 8248 5457 8276
rect 5399 8245 5411 8248
rect 5353 8239 5411 8245
rect 5445 8245 5457 8248
rect 5491 8276 5503 8279
rect 6270 8276 6276 8288
rect 5491 8248 6276 8276
rect 5491 8245 5503 8248
rect 5445 8239 5503 8245
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 12710 8276 12716 8288
rect 7892 8248 12716 8276
rect 7892 8236 7898 8248
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 13004 8276 13032 8384
rect 13538 8372 13544 8424
rect 13596 8372 13602 8424
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 14844 8412 14872 8452
rect 15654 8440 15660 8492
rect 15712 8440 15718 8492
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16172 8452 17233 8480
rect 16172 8440 16178 8452
rect 17221 8449 17233 8452
rect 17267 8480 17279 8483
rect 17310 8480 17316 8492
rect 17267 8452 17316 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 17586 8480 17592 8492
rect 17512 8452 17592 8480
rect 13771 8384 14872 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 14918 8372 14924 8424
rect 14976 8372 14982 8424
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 15620 8384 16681 8412
rect 15620 8372 15626 8384
rect 16669 8381 16681 8384
rect 16715 8412 16727 8415
rect 16758 8412 16764 8424
rect 16715 8384 16764 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 17512 8412 17540 8452
rect 17586 8440 17592 8452
rect 17644 8480 17650 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17644 8452 18613 8480
rect 17644 8440 17650 8452
rect 18601 8449 18613 8452
rect 18647 8480 18659 8483
rect 18874 8480 18880 8492
rect 18647 8452 18880 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 16908 8384 17540 8412
rect 16908 8372 16914 8384
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 19426 8412 19432 8424
rect 18748 8384 19432 8412
rect 18748 8372 18754 8384
rect 19426 8372 19432 8384
rect 19484 8372 19490 8424
rect 13081 8347 13139 8353
rect 13081 8313 13093 8347
rect 13127 8344 13139 8347
rect 13906 8344 13912 8356
rect 13127 8316 13912 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 19576 8316 22094 8344
rect 19576 8304 19582 8316
rect 16850 8276 16856 8288
rect 13004 8248 16856 8276
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 22066 8276 22094 8316
rect 23658 8276 23664 8288
rect 22066 8248 23664 8276
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2130 8072 2136 8084
rect 1627 8044 2136 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 2556 8044 5365 8072
rect 2556 8032 2562 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7558 8072 7564 8084
rect 7064 8044 7564 8072
rect 7064 8032 7070 8044
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 8570 8032 8576 8084
rect 8628 8032 8634 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 9732 8044 11161 8072
rect 9732 8032 9738 8044
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 11149 8035 11207 8041
rect 12342 8032 12348 8084
rect 12400 8032 12406 8084
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13630 8072 13636 8084
rect 13495 8044 13636 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14734 8072 14740 8084
rect 14323 8044 14740 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 16761 8075 16819 8081
rect 16761 8072 16773 8075
rect 14884 8044 16773 8072
rect 14884 8032 14890 8044
rect 16761 8041 16773 8044
rect 16807 8041 16819 8075
rect 16761 8035 16819 8041
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 18785 8075 18843 8081
rect 18785 8072 18797 8075
rect 17460 8044 18797 8072
rect 17460 8032 17466 8044
rect 18785 8041 18797 8044
rect 18831 8041 18843 8075
rect 18785 8035 18843 8041
rect 750 7964 756 8016
rect 808 8004 814 8016
rect 3973 8007 4031 8013
rect 808 7976 2774 8004
rect 808 7964 814 7976
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2406 7936 2412 7948
rect 2271 7908 2412 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1360 7840 1777 7868
rect 1360 7828 1366 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 2746 7868 2774 7976
rect 3973 7973 3985 8007
rect 4019 8004 4031 8007
rect 7650 8004 7656 8016
rect 4019 7976 7656 8004
rect 4019 7973 4031 7976
rect 3973 7967 4031 7973
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 9858 8004 9864 8016
rect 7944 7976 9864 8004
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 5718 7936 5724 7948
rect 2915 7908 5724 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 2746 7840 4169 7868
rect 1765 7831 1823 7837
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 1780 7732 1808 7831
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 5592 7840 5917 7868
rect 5592 7828 5598 7840
rect 5905 7837 5917 7840
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6178 7828 6184 7880
rect 6236 7828 6242 7880
rect 7944 7877 7972 7976
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 7973 10195 8007
rect 10137 7967 10195 7973
rect 9398 7896 9404 7948
rect 9456 7896 9462 7948
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9858 7868 9864 7880
rect 9324 7840 9864 7868
rect 3513 7803 3571 7809
rect 3513 7800 3525 7803
rect 2746 7772 3525 7800
rect 2746 7732 2774 7772
rect 3513 7769 3525 7772
rect 3559 7769 3571 7803
rect 6730 7800 6736 7812
rect 3513 7763 3571 7769
rect 4724 7772 6736 7800
rect 1780 7704 2774 7732
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 4724 7741 4752 7772
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 7466 7760 7472 7812
rect 7524 7800 7530 7812
rect 9324 7800 9352 7840
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 7524 7772 9352 7800
rect 10152 7800 10180 7967
rect 11330 7964 11336 8016
rect 11388 8004 11394 8016
rect 17221 8007 17279 8013
rect 17221 8004 17233 8007
rect 11388 7976 17233 8004
rect 11388 7964 11394 7976
rect 17221 7973 17233 7976
rect 17267 7973 17279 8007
rect 17221 7967 17279 7973
rect 10594 7896 10600 7948
rect 10652 7896 10658 7948
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 10827 7908 12664 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7868 10563 7871
rect 10686 7868 10692 7880
rect 10551 7840 10692 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11296 7840 11713 7868
rect 11296 7828 11302 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 12434 7800 12440 7812
rect 10152 7772 12440 7800
rect 7524 7760 7530 7772
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 12636 7800 12664 7908
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 14737 7939 14795 7945
rect 14737 7936 14749 7939
rect 12768 7908 14749 7936
rect 12768 7896 12774 7908
rect 14737 7905 14749 7908
rect 14783 7905 14795 7939
rect 14737 7899 14795 7905
rect 14921 7939 14979 7945
rect 14921 7905 14933 7939
rect 14967 7936 14979 7939
rect 17126 7936 17132 7948
rect 14967 7908 17132 7936
rect 14967 7905 14979 7908
rect 14921 7899 14979 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 13446 7868 13452 7880
rect 12851 7840 13452 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 14240 7840 15485 7868
rect 14240 7828 14246 7840
rect 15473 7837 15485 7840
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 16022 7828 16028 7880
rect 16080 7868 16086 7880
rect 16117 7871 16175 7877
rect 16117 7868 16129 7871
rect 16080 7840 16129 7868
rect 16080 7828 16086 7840
rect 16117 7837 16129 7840
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 15286 7800 15292 7812
rect 12636 7772 15292 7800
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 16132 7800 16160 7831
rect 16206 7828 16212 7880
rect 16264 7868 16270 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 16264 7840 17417 7868
rect 16264 7828 16270 7840
rect 17405 7837 17417 7840
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18414 7868 18420 7880
rect 18187 7840 18420 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 17770 7800 17776 7812
rect 16132 7772 17776 7800
rect 17770 7760 17776 7772
rect 17828 7760 17834 7812
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 3292 7704 3341 7732
rect 3292 7692 3298 7704
rect 3329 7701 3341 7704
rect 3375 7701 3387 7735
rect 3329 7695 3387 7701
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7701 4767 7735
rect 4709 7695 4767 7701
rect 5626 7692 5632 7744
rect 5684 7692 5690 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7374 7732 7380 7744
rect 6972 7704 7380 7732
rect 6972 7692 6978 7704
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 8720 7704 9873 7732
rect 8720 7692 8726 7704
rect 9861 7701 9873 7704
rect 9907 7732 9919 7735
rect 10042 7732 10048 7744
rect 9907 7704 10048 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 10042 7692 10048 7704
rect 10100 7732 10106 7744
rect 11054 7732 11060 7744
rect 10100 7704 11060 7732
rect 10100 7692 10106 7704
rect 11054 7692 11060 7704
rect 11112 7732 11118 7744
rect 11333 7735 11391 7741
rect 11333 7732 11345 7735
rect 11112 7704 11345 7732
rect 11112 7692 11118 7704
rect 11333 7701 11345 7704
rect 11379 7701 11391 7735
rect 11333 7695 11391 7701
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 4522 7488 4528 7540
rect 4580 7488 4586 7540
rect 4706 7488 4712 7540
rect 4764 7488 4770 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5350 7528 5356 7540
rect 4939 7500 5356 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 7101 7531 7159 7537
rect 7101 7528 7113 7531
rect 6328 7500 7113 7528
rect 6328 7488 6334 7500
rect 7101 7497 7113 7500
rect 7147 7528 7159 7531
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 7147 7500 7941 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 10778 7528 10784 7540
rect 9631 7500 10784 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11241 7531 11299 7537
rect 11241 7528 11253 7531
rect 11112 7500 11253 7528
rect 11112 7488 11118 7500
rect 11241 7497 11253 7500
rect 11287 7497 11299 7531
rect 11241 7491 11299 7497
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12066 7528 12072 7540
rect 11839 7500 12072 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 13722 7488 13728 7540
rect 13780 7488 13786 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15252 7500 16037 7528
rect 15252 7488 15258 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 24026 7488 24032 7540
rect 24084 7488 24090 7540
rect 3620 7432 15056 7460
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2222 7392 2228 7404
rect 1903 7364 2228 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 3620 7401 3648 7432
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6270 7392 6276 7404
rect 6043 7364 6276 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 7098 7392 7104 7404
rect 6687 7364 7104 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7834 7392 7840 7404
rect 7524 7364 7840 7392
rect 7524 7352 7530 7364
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8662 7392 8668 7404
rect 8343 7364 8668 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8938 7352 8944 7404
rect 8996 7392 9002 7404
rect 10502 7392 10508 7404
rect 8996 7364 10508 7392
rect 8996 7352 9002 7364
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12342 7392 12348 7404
rect 12023 7364 12348 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13354 7392 13360 7404
rect 13127 7364 13360 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13872 7364 14289 7392
rect 13872 7352 13878 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 2866 7324 2872 7336
rect 1627 7296 2872 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 2866 7284 2872 7296
rect 2924 7284 2930 7336
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4706 7324 4712 7336
rect 3375 7296 4712 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 5626 7324 5632 7336
rect 5215 7296 5632 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 6972 7296 8585 7324
rect 6972 7284 6978 7296
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8754 7284 8760 7336
rect 8812 7324 8818 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 8812 7296 10701 7324
rect 8812 7284 8818 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 6178 7256 6184 7268
rect 2746 7228 6184 7256
rect 658 7148 664 7200
rect 716 7188 722 7200
rect 2746 7188 2774 7228
rect 6178 7216 6184 7228
rect 6236 7216 6242 7268
rect 7469 7259 7527 7265
rect 7469 7256 7481 7259
rect 7300 7228 7481 7256
rect 716 7160 2774 7188
rect 716 7148 722 7160
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7300 7188 7328 7228
rect 7469 7225 7481 7228
rect 7515 7225 7527 7259
rect 7469 7219 7527 7225
rect 10226 7216 10232 7268
rect 10284 7216 10290 7268
rect 10888 7256 10916 7287
rect 11514 7284 11520 7336
rect 11572 7324 11578 7336
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 11572 7296 14933 7324
rect 11572 7284 11578 7296
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 15028 7324 15056 7432
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 15160 7432 16865 7460
rect 15160 7420 15166 7432
rect 16853 7429 16865 7432
rect 16899 7429 16911 7463
rect 16853 7423 16911 7429
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 20680 7364 22293 7392
rect 20680 7352 20686 7364
rect 22281 7361 22293 7364
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 23658 7352 23664 7404
rect 23716 7392 23722 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 23716 7364 24317 7392
rect 23716 7352 23722 7364
rect 24305 7361 24317 7364
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 21082 7324 21088 7336
rect 15028 7296 21088 7324
rect 14921 7287 14979 7293
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 16022 7256 16028 7268
rect 10888 7228 16028 7256
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 7064 7160 7328 7188
rect 7745 7191 7803 7197
rect 7064 7148 7070 7160
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 7834 7188 7840 7200
rect 7791 7160 7840 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 7834 7148 7840 7160
rect 7892 7188 7898 7200
rect 12158 7188 12164 7200
rect 7892 7160 12164 7188
rect 7892 7148 7898 7160
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12342 7148 12348 7200
rect 12400 7148 12406 7200
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 13354 7188 13360 7200
rect 12575 7160 13360 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 6822 6984 6828 6996
rect 2746 6956 6828 6984
rect 106 6876 112 6928
rect 164 6916 170 6928
rect 2746 6916 2774 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7190 6944 7196 6996
rect 7248 6944 7254 6996
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7834 6984 7840 6996
rect 7432 6956 7840 6984
rect 7432 6944 7438 6956
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 164 6888 2774 6916
rect 164 6876 170 6888
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 15930 6916 15936 6928
rect 5684 6888 15936 6916
rect 5684 6876 5690 6888
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 1946 6848 1952 6860
rect 1903 6820 1952 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2866 6848 2872 6860
rect 2731 6820 2872 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3973 6851 4031 6857
rect 3292 6820 3832 6848
rect 3292 6808 3298 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 2774 6780 2780 6792
rect 1627 6752 2780 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3694 6780 3700 6792
rect 2832 6752 3700 6780
rect 2832 6740 2838 6752
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 3804 6780 3832 6820
rect 3973 6817 3985 6851
rect 4019 6848 4031 6851
rect 4154 6848 4160 6860
rect 4019 6820 4160 6848
rect 4019 6817 4031 6820
rect 3973 6811 4031 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4264 6820 5948 6848
rect 4264 6780 4292 6820
rect 3804 6752 4292 6780
rect 4893 6783 4951 6789
rect 4893 6749 4905 6783
rect 4939 6780 4951 6783
rect 5350 6780 5356 6792
rect 4939 6752 5356 6780
rect 4939 6749 4951 6752
rect 4893 6743 4951 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 3329 6715 3387 6721
rect 3329 6712 3341 6715
rect 1360 6684 3341 6712
rect 1360 6672 1366 6684
rect 3329 6681 3341 6684
rect 3375 6681 3387 6715
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 3329 6675 3387 6681
rect 3712 6684 4169 6712
rect 474 6604 480 6656
rect 532 6644 538 6656
rect 3712 6644 3740 6684
rect 4157 6681 4169 6684
rect 4203 6712 4215 6715
rect 4249 6715 4307 6721
rect 4249 6712 4261 6715
rect 4203 6684 4261 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 4249 6681 4261 6684
rect 4295 6681 4307 6715
rect 4249 6675 4307 6681
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5920 6712 5948 6820
rect 7650 6808 7656 6860
rect 7708 6808 7714 6860
rect 10318 6808 10324 6860
rect 10376 6808 10382 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 11940 6820 12173 6848
rect 11940 6808 11946 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 21361 6851 21419 6857
rect 12161 6811 12219 6817
rect 12406 6820 15148 6848
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7892 6752 7941 6780
rect 7892 6740 7898 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 7377 6715 7435 6721
rect 5132 6684 5856 6712
rect 5920 6684 7236 6712
rect 5132 6672 5138 6684
rect 532 6616 3740 6644
rect 5169 6647 5227 6653
rect 532 6604 538 6616
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5534 6644 5540 6656
rect 5215 6616 5540 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5828 6653 5856 6684
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6613 5871 6647
rect 5813 6607 5871 6613
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6914 6644 6920 6656
rect 6503 6616 6920 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 7098 6644 7104 6656
rect 7055 6616 7104 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7208 6644 7236 6684
rect 7377 6681 7389 6715
rect 7423 6712 7435 6715
rect 8478 6712 8484 6724
rect 7423 6684 8484 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 9140 6712 9168 6743
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11606 6780 11612 6792
rect 11563 6752 11612 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 12406 6780 12434 6820
rect 11848 6752 12434 6780
rect 11848 6740 11854 6752
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 15120 6789 15148 6820
rect 21361 6817 21373 6851
rect 21407 6848 21419 6851
rect 22554 6848 22560 6860
rect 21407 6820 22560 6848
rect 21407 6817 21419 6820
rect 21361 6811 21419 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 20714 6740 20720 6792
rect 20772 6740 20778 6792
rect 10502 6712 10508 6724
rect 9140 6684 10508 6712
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 10870 6672 10876 6724
rect 10928 6672 10934 6724
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6681 11115 6715
rect 11057 6675 11115 6681
rect 10778 6644 10784 6656
rect 7208 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11072 6644 11100 6675
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12400 6684 13277 6712
rect 12400 6672 12406 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 14090 6644 14096 6656
rect 11072 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14921 6647 14979 6653
rect 14921 6613 14933 6647
rect 14967 6644 14979 6647
rect 18506 6644 18512 6656
rect 14967 6616 18512 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 18506 6604 18512 6616
rect 18564 6604 18570 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6440 3111 6443
rect 3602 6440 3608 6452
rect 3099 6412 3608 6440
rect 3099 6409 3111 6412
rect 3053 6403 3111 6409
rect 3234 6372 3240 6384
rect 1872 6344 3240 6372
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1872 6313 1900 6344
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3528 6313 3556 6412
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4062 6440 4068 6452
rect 4019 6412 4068 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 5994 6440 6000 6452
rect 5859 6412 6000 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6822 6440 6828 6452
rect 6227 6412 6828 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 9585 6443 9643 6449
rect 9585 6409 9597 6443
rect 9631 6440 9643 6443
rect 10594 6440 10600 6452
rect 9631 6412 10600 6440
rect 9631 6409 9643 6412
rect 9585 6403 9643 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 11480 6412 12173 6440
rect 11480 6400 11486 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14642 6440 14648 6452
rect 14323 6412 14648 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 21910 6372 21916 6384
rect 5408 6344 21916 6372
rect 5408 6332 5414 6344
rect 21910 6332 21916 6344
rect 21968 6332 21974 6384
rect 23937 6375 23995 6381
rect 23937 6341 23949 6375
rect 23983 6372 23995 6375
rect 28718 6372 28724 6384
rect 23983 6344 28724 6372
rect 23983 6341 23995 6344
rect 23937 6335 23995 6341
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 4396 6276 5457 6304
rect 4396 6264 4402 6276
rect 5445 6273 5457 6276
rect 5491 6304 5503 6307
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 5491 6276 5917 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 9398 6304 9404 6316
rect 5905 6267 5963 6273
rect 6104 6276 9404 6304
rect 566 6196 572 6248
rect 624 6236 630 6248
rect 6104 6236 6132 6276
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 9548 6276 10333 6304
rect 9548 6264 9554 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10468 6276 10885 6304
rect 10468 6264 10474 6276
rect 10873 6273 10885 6276
rect 10919 6304 10931 6307
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10919 6276 10977 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12342 6304 12348 6316
rect 11756 6276 12348 6304
rect 11756 6264 11762 6276
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12802 6264 12808 6316
rect 12860 6304 12866 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12860 6276 12909 6304
rect 12860 6264 12866 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 22278 6264 22284 6316
rect 22336 6304 22342 6316
rect 23017 6307 23075 6313
rect 23017 6304 23029 6307
rect 22336 6276 23029 6304
rect 22336 6264 22342 6276
rect 23017 6273 23029 6276
rect 23063 6304 23075 6307
rect 23952 6304 23980 6335
rect 28718 6332 28724 6344
rect 28776 6332 28782 6384
rect 23063 6276 23980 6304
rect 23063 6273 23075 6276
rect 23017 6267 23075 6273
rect 624 6208 6132 6236
rect 624 6196 630 6208
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6696 6208 6929 6236
rect 6696 6196 6702 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8895 6208 8953 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 8941 6205 8953 6208
rect 8987 6236 8999 6239
rect 9674 6236 9680 6248
rect 8987 6208 9680 6236
rect 8987 6205 8999 6208
rect 8941 6199 8999 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 12032 6208 13553 6236
rect 12032 6196 12038 6208
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 4430 6168 4436 6180
rect 3375 6140 4436 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 13998 6168 14004 6180
rect 7064 6140 14004 6168
rect 7064 6128 7070 6140
rect 13998 6128 14004 6140
rect 14056 6128 14062 6180
rect 24026 6168 24032 6180
rect 23308 6140 24032 6168
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 4154 6100 4160 6112
rect 1912 6072 4160 6100
rect 1912 6060 1918 6072
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 6914 6100 6920 6112
rect 5307 6072 6920 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 16666 6100 16672 6112
rect 7156 6072 16672 6100
rect 7156 6060 7162 6072
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 23308 6109 23336 6140
rect 24026 6128 24032 6140
rect 24084 6128 24090 6180
rect 23293 6103 23351 6109
rect 23293 6069 23305 6103
rect 23339 6069 23351 6103
rect 23293 6063 23351 6069
rect 23477 6103 23535 6109
rect 23477 6069 23489 6103
rect 23523 6100 23535 6103
rect 23566 6100 23572 6112
rect 23523 6072 23572 6100
rect 23523 6069 23535 6072
rect 23477 6063 23535 6069
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2556 5868 2881 5896
rect 2556 5856 2562 5868
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 5261 5899 5319 5905
rect 5261 5865 5273 5899
rect 5307 5896 5319 5899
rect 9030 5896 9036 5908
rect 5307 5868 9036 5896
rect 5307 5865 5319 5868
rect 5261 5859 5319 5865
rect 3988 5828 4016 5859
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9306 5896 9312 5908
rect 9171 5868 9312 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9766 5896 9772 5908
rect 9723 5868 9772 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 11701 5899 11759 5905
rect 11701 5865 11713 5899
rect 11747 5896 11759 5899
rect 16850 5896 16856 5908
rect 11747 5868 16856 5896
rect 11747 5865 11759 5868
rect 11701 5859 11759 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19518 5896 19524 5908
rect 19383 5868 19524 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 22833 5899 22891 5905
rect 22833 5865 22845 5899
rect 22879 5896 22891 5899
rect 26234 5896 26240 5908
rect 22879 5868 26240 5896
rect 22879 5865 22891 5868
rect 22833 5859 22891 5865
rect 6362 5828 6368 5840
rect 3988 5800 6368 5828
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 7800 5800 12434 5828
rect 7800 5788 7806 5800
rect 1854 5720 1860 5772
rect 1912 5720 1918 5772
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 2746 5732 3341 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2746 5692 2774 5732
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 3510 5760 3516 5772
rect 3375 5732 3516 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 4028 5732 5733 5760
rect 4028 5720 4034 5732
rect 1627 5664 2774 5692
rect 3053 5695 3111 5701
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5692 3663 5695
rect 4154 5692 4160 5704
rect 3651 5664 4160 5692
rect 3651 5661 3663 5664
rect 3605 5655 3663 5661
rect 3068 5624 3096 5655
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4614 5692 4620 5704
rect 4264 5664 4620 5692
rect 3510 5624 3516 5636
rect 3068 5596 3516 5624
rect 3510 5584 3516 5596
rect 3568 5624 3574 5636
rect 3878 5624 3884 5636
rect 3568 5596 3884 5624
rect 3568 5584 3574 5596
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 4264 5556 4292 5664
rect 4614 5652 4620 5664
rect 4672 5692 4678 5704
rect 5460 5701 5488 5732
rect 5721 5729 5733 5732
rect 5767 5729 5779 5763
rect 5721 5723 5779 5729
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 6604 5732 11928 5760
rect 6604 5720 6610 5732
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4672 5664 4813 5692
rect 4672 5652 4678 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 11900 5701 11928 5732
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 9180 5664 9321 5692
rect 9180 5652 9186 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5661 11943 5695
rect 12406 5692 12434 5800
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 14550 5760 14556 5772
rect 13780 5732 14556 5760
rect 13780 5720 13786 5732
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 14829 5763 14887 5769
rect 14829 5760 14841 5763
rect 14792 5732 14841 5760
rect 14792 5720 14798 5732
rect 14829 5729 14841 5732
rect 14875 5729 14887 5763
rect 14829 5723 14887 5729
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 17092 5732 17141 5760
rect 17092 5720 17098 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 18877 5763 18935 5769
rect 18877 5729 18889 5763
rect 18923 5760 18935 5763
rect 20714 5760 20720 5772
rect 18923 5732 20720 5760
rect 18923 5729 18935 5732
rect 18877 5723 18935 5729
rect 20714 5720 20720 5732
rect 20772 5720 20778 5772
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 12406 5664 13645 5692
rect 11885 5655 11943 5661
rect 13633 5661 13645 5664
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 22332 5695 22390 5701
rect 22332 5692 22344 5695
rect 14369 5655 14427 5661
rect 22066 5664 22344 5692
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 14384 5624 14412 5655
rect 6788 5596 14412 5624
rect 6788 5584 6794 5596
rect 14550 5584 14556 5636
rect 14608 5624 14614 5636
rect 14608 5596 15332 5624
rect 14608 5584 14614 5596
rect 2372 5528 4292 5556
rect 4617 5559 4675 5565
rect 2372 5516 2378 5528
rect 4617 5525 4629 5559
rect 4663 5556 4675 5559
rect 6454 5556 6460 5568
rect 4663 5528 6460 5556
rect 4663 5525 4675 5528
rect 4617 5519 4675 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 10744 5528 12817 5556
rect 10744 5516 10750 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 12805 5519 12863 5525
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 15102 5556 15108 5568
rect 13495 5528 15108 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 15304 5556 15332 5596
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 16356 5596 17417 5624
rect 16356 5584 16362 5596
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 19426 5624 19432 5636
rect 18630 5596 19432 5624
rect 17405 5587 17463 5593
rect 19426 5584 19432 5596
rect 19484 5584 19490 5636
rect 16577 5559 16635 5565
rect 16577 5556 16589 5559
rect 15304 5528 16589 5556
rect 16577 5525 16589 5528
rect 16623 5556 16635 5559
rect 22066 5556 22094 5664
rect 22332 5661 22344 5664
rect 22378 5692 22390 5695
rect 22848 5692 22876 5859
rect 26234 5856 26240 5868
rect 26292 5856 26298 5908
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 25961 5763 26019 5769
rect 25961 5760 25973 5763
rect 23532 5732 25973 5760
rect 23532 5720 23538 5732
rect 25961 5729 25973 5732
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 26694 5720 26700 5772
rect 26752 5720 26758 5772
rect 22378 5664 22876 5692
rect 25777 5695 25835 5701
rect 22378 5661 22390 5664
rect 22332 5655 22390 5661
rect 25777 5661 25789 5695
rect 25823 5661 25835 5695
rect 25777 5655 25835 5661
rect 22419 5627 22477 5633
rect 22419 5593 22431 5627
rect 22465 5624 22477 5627
rect 24762 5624 24768 5636
rect 22465 5596 24768 5624
rect 22465 5593 22477 5596
rect 22419 5587 22477 5593
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 25792 5624 25820 5655
rect 27522 5624 27528 5636
rect 25792 5596 27528 5624
rect 27522 5584 27528 5596
rect 27580 5584 27586 5636
rect 16623 5528 22094 5556
rect 16623 5525 16635 5528
rect 16577 5519 16635 5525
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 4062 5352 4068 5364
rect 1872 5324 4068 5352
rect 1872 5225 1900 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 5718 5352 5724 5364
rect 4203 5324 5724 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 22278 5352 22284 5364
rect 21836 5324 22284 5352
rect 3786 5284 3792 5296
rect 3068 5256 3792 5284
rect 3068 5225 3096 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 4430 5284 4436 5296
rect 3896 5256 4436 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 3896 5216 3924 5256
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 4893 5287 4951 5293
rect 4893 5284 4905 5287
rect 4540 5256 4905 5284
rect 4540 5228 4568 5256
rect 4893 5253 4905 5256
rect 4939 5253 4951 5287
rect 4893 5247 4951 5253
rect 3743 5188 3924 5216
rect 4341 5219 4399 5225
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4522 5216 4528 5228
rect 4387 5188 4528 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4614 5176 4620 5228
rect 4672 5176 4678 5228
rect 20898 5176 20904 5228
rect 20956 5216 20962 5228
rect 21836 5225 21864 5324
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22419 5355 22477 5361
rect 22419 5321 22431 5355
rect 22465 5352 22477 5355
rect 23474 5352 23480 5364
rect 22465 5324 23480 5352
rect 22465 5321 22477 5324
rect 22419 5315 22477 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 24762 5244 24768 5296
rect 24820 5284 24826 5296
rect 24949 5287 25007 5293
rect 24949 5284 24961 5287
rect 24820 5256 24961 5284
rect 24820 5244 24826 5256
rect 24949 5253 24961 5256
rect 24995 5253 25007 5287
rect 24949 5247 25007 5253
rect 26605 5287 26663 5293
rect 26605 5253 26617 5287
rect 26651 5284 26663 5287
rect 27614 5284 27620 5296
rect 26651 5256 27620 5284
rect 26651 5253 26663 5256
rect 26605 5247 26663 5253
rect 27614 5244 27620 5256
rect 27672 5284 27678 5296
rect 28534 5284 28540 5296
rect 27672 5256 28540 5284
rect 27672 5244 27678 5256
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 28997 5287 29055 5293
rect 28997 5253 29009 5287
rect 29043 5284 29055 5287
rect 29086 5284 29092 5296
rect 29043 5256 29092 5284
rect 29043 5253 29055 5256
rect 28997 5247 29055 5253
rect 29086 5244 29092 5256
rect 29144 5244 29150 5296
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 20956 5188 21833 5216
rect 20956 5176 20962 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22348 5219 22406 5225
rect 22348 5185 22360 5219
rect 22394 5216 22406 5219
rect 23566 5216 23572 5228
rect 22394 5188 23572 5216
rect 22394 5185 22406 5188
rect 22348 5179 22406 5185
rect 23566 5176 23572 5188
rect 23624 5176 23630 5228
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 1636 5120 4997 5148
rect 1636 5108 1642 5120
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 24765 5151 24823 5157
rect 24765 5117 24777 5151
rect 24811 5117 24823 5151
rect 24765 5111 24823 5117
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5117 27215 5151
rect 27157 5111 27215 5117
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5080 3571 5083
rect 6086 5080 6092 5092
rect 3559 5052 6092 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 18598 5040 18604 5092
rect 18656 5080 18662 5092
rect 21358 5080 21364 5092
rect 18656 5052 21364 5080
rect 18656 5040 18662 5052
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 24780 5080 24808 5111
rect 25498 5080 25504 5092
rect 24780 5052 25504 5080
rect 25498 5040 25504 5052
rect 25556 5040 25562 5092
rect 27172 5080 27200 5111
rect 27338 5108 27344 5160
rect 27396 5108 27402 5160
rect 29457 5151 29515 5157
rect 29457 5117 29469 5151
rect 29503 5117 29515 5151
rect 29457 5111 29515 5117
rect 29086 5080 29092 5092
rect 27172 5052 29092 5080
rect 29086 5040 29092 5052
rect 29144 5040 29150 5092
rect 29472 5080 29500 5111
rect 29638 5108 29644 5160
rect 29696 5108 29702 5160
rect 31297 5151 31355 5157
rect 31297 5117 31309 5151
rect 31343 5148 31355 5151
rect 31754 5148 31760 5160
rect 31343 5120 31760 5148
rect 31343 5117 31355 5120
rect 31297 5111 31355 5117
rect 31754 5108 31760 5120
rect 31812 5148 31818 5160
rect 32490 5148 32496 5160
rect 31812 5120 32496 5148
rect 31812 5108 31818 5120
rect 32490 5108 32496 5120
rect 32548 5108 32554 5160
rect 32858 5080 32864 5092
rect 29472 5052 32864 5080
rect 32858 5040 32864 5052
rect 32916 5040 32922 5092
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 4982 5012 4988 5024
rect 2915 4984 4988 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20772 4984 21005 5012
rect 20772 4972 20778 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3326 4808 3332 4820
rect 2915 4780 3332 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3421 4811 3479 4817
rect 3421 4777 3433 4811
rect 3467 4808 3479 4811
rect 3510 4808 3516 4820
rect 3467 4780 3516 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3786 4808 3792 4820
rect 3651 4780 3792 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 10134 4808 10140 4820
rect 4120 4780 10140 4808
rect 4120 4768 4126 4780
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 14921 4811 14979 4817
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 16298 4808 16304 4820
rect 14967 4780 16304 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 19521 4811 19579 4817
rect 19521 4777 19533 4811
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 23063 4811 23121 4817
rect 23063 4777 23075 4811
rect 23109 4808 23121 4811
rect 27338 4808 27344 4820
rect 23109 4780 27344 4808
rect 23109 4777 23121 4780
rect 23063 4771 23121 4777
rect 3973 4743 4031 4749
rect 3973 4709 3985 4743
rect 4019 4740 4031 4743
rect 9950 4740 9956 4752
rect 4019 4712 9956 4740
rect 4019 4709 4031 4712
rect 3973 4703 4031 4709
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 19536 4740 19564 4771
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 14292 4712 19564 4740
rect 24719 4743 24777 4749
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 1360 4644 1593 4672
rect 1360 4632 1366 4644
rect 1581 4641 1593 4644
rect 1627 4672 1639 4675
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 1627 4644 4629 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 4617 4635 4675 4641
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4764 4644 4813 4672
rect 4764 4632 4770 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 1857 4607 1915 4613
rect 1857 4573 1869 4607
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 1872 4536 1900 4567
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2648 4576 3065 4604
rect 2648 4564 2654 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3418 4604 3424 4616
rect 3099 4576 3424 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4246 4604 4252 4616
rect 4203 4576 4252 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4246 4564 4252 4576
rect 4304 4604 4310 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4304 4576 4445 4604
rect 4304 4564 4310 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 14292 4613 14320 4712
rect 24719 4709 24731 4743
rect 24765 4740 24777 4743
rect 29638 4740 29644 4752
rect 24765 4712 29644 4740
rect 24765 4709 24777 4712
rect 24719 4703 24777 4709
rect 29638 4700 29644 4712
rect 29696 4700 29702 4752
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15160 4644 15761 4672
rect 15160 4632 15166 4644
rect 15749 4641 15761 4644
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 17402 4632 17408 4684
rect 17460 4632 17466 4684
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 19944 4644 23336 4672
rect 19944 4632 19950 4644
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 11112 4576 14289 4604
rect 11112 4564 11118 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 19475 4576 20269 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20257 4573 20269 4576
rect 20303 4604 20315 4607
rect 20898 4604 20904 4616
rect 20303 4576 20904 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21358 4564 21364 4616
rect 21416 4604 21422 4616
rect 22960 4607 23018 4613
rect 22960 4604 22972 4607
rect 21416 4576 22972 4604
rect 21416 4564 21422 4576
rect 22960 4573 22972 4576
rect 23006 4573 23018 4607
rect 23308 4604 23336 4644
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 23308 4576 24628 4604
rect 22960 4567 23018 4573
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 8846 4536 8852 4548
rect 1872 4508 8852 4536
rect 8846 4496 8852 4508
rect 8904 4496 8910 4548
rect 13814 4496 13820 4548
rect 13872 4536 13878 4548
rect 15933 4539 15991 4545
rect 15933 4536 15945 4539
rect 13872 4508 15945 4536
rect 13872 4496 13878 4508
rect 15933 4505 15945 4508
rect 15979 4536 15991 4539
rect 23566 4536 23572 4548
rect 15979 4508 23572 4536
rect 15979 4505 15991 4508
rect 15933 4499 15991 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 19886 4428 19892 4480
rect 19944 4428 19950 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2038 4128 2044 4140
rect 1903 4100 2044 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2832 4100 3065 4128
rect 2832 4088 2838 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3752 4100 3985 4128
rect 3752 4088 3758 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 16850 4088 16856 4140
rect 16908 4088 16914 4140
rect 1596 4060 1624 4088
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 1596 4032 4169 4060
rect 4157 4029 4169 4032
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 14148 4032 17049 4060
rect 14148 4020 14154 4032
rect 17037 4029 17049 4032
rect 17083 4060 17095 4063
rect 18598 4060 18604 4072
rect 17083 4032 18604 4060
rect 17083 4029 17095 4032
rect 17037 4023 17095 4029
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4060 18751 4063
rect 20070 4060 20076 4072
rect 18739 4032 20076 4060
rect 18739 4029 18751 4032
rect 18693 4023 18751 4029
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 382 3952 388 4004
rect 440 3992 446 4004
rect 2869 3995 2927 4001
rect 2869 3992 2881 3995
rect 440 3964 2881 3992
rect 440 3952 446 3964
rect 2869 3961 2881 3964
rect 2915 3961 2927 3995
rect 2869 3955 2927 3961
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 8938 3992 8944 4004
rect 3559 3964 8944 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 8938 3952 8944 3964
rect 8996 3952 9002 4004
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 2832 3692 3525 3720
rect 2832 3680 2838 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 3513 3683 3571 3689
rect 3973 3723 4031 3729
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 7558 3720 7564 3732
rect 4019 3692 7564 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 12434 3720 12440 3732
rect 12207 3692 12440 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 12434 3680 12440 3692
rect 12492 3720 12498 3732
rect 13722 3720 13728 3732
rect 12492 3692 13728 3720
rect 12492 3680 12498 3692
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 32490 3680 32496 3732
rect 32548 3720 32554 3732
rect 41414 3720 41420 3732
rect 32548 3692 41420 3720
rect 32548 3680 32554 3692
rect 41414 3680 41420 3692
rect 41472 3680 41478 3732
rect 2866 3612 2872 3664
rect 2924 3612 2930 3664
rect 3418 3612 3424 3664
rect 3476 3612 3482 3664
rect 29178 3612 29184 3664
rect 29236 3652 29242 3664
rect 44082 3652 44088 3664
rect 29236 3624 44088 3652
rect 29236 3612 29242 3624
rect 44082 3612 44088 3624
rect 44140 3612 44146 3664
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 1360 3556 1593 3584
rect 1360 3544 1366 3556
rect 1581 3553 1593 3556
rect 1627 3584 1639 3587
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 1627 3556 4629 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 26694 3544 26700 3596
rect 26752 3584 26758 3596
rect 46750 3584 46756 3596
rect 26752 3556 46756 3584
rect 26752 3544 26758 3556
rect 46750 3544 46756 3556
rect 46808 3544 46814 3596
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3326 3516 3332 3528
rect 3099 3488 3332 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 1872 3448 1900 3479
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4120 3488 4169 3516
rect 4120 3476 4126 3488
rect 4157 3485 4169 3488
rect 4203 3516 4215 3519
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4203 3488 4445 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 49418 3516 49424 3528
rect 27672 3488 49424 3516
rect 27672 3476 27678 3488
rect 49418 3476 49424 3488
rect 49476 3476 49482 3528
rect 7466 3448 7472 3460
rect 1872 3420 7472 3448
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 38746 3448 38752 3460
rect 19392 3420 38752 3448
rect 19392 3408 19398 3420
rect 38746 3408 38752 3420
rect 38804 3408 38810 3460
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3234 3176 3240 3188
rect 2915 3148 3240 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 3559 3148 7144 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 1210 3068 1216 3120
rect 1268 3108 1274 3120
rect 7116 3108 7144 3148
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 10597 3179 10655 3185
rect 8352 3148 10456 3176
rect 8352 3136 8358 3148
rect 8754 3108 8760 3120
rect 1268 3080 3740 3108
rect 7116 3080 8760 3108
rect 1268 3068 1274 3080
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3712 3049 3740 3080
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 10428 3108 10456 3148
rect 10597 3145 10609 3179
rect 10643 3176 10655 3179
rect 11054 3176 11060 3188
rect 10643 3148 11060 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 11164 3148 12725 3176
rect 11164 3108 11192 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 12713 3139 12771 3145
rect 10428 3080 11192 3108
rect 11793 3111 11851 3117
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 12434 3108 12440 3120
rect 11839 3080 12440 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3108 12679 3111
rect 13814 3108 13820 3120
rect 12667 3080 13820 3108
rect 12667 3077 12679 3080
rect 12621 3071 12679 3077
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 14090 3068 14096 3120
rect 14148 3068 14154 3120
rect 15841 3111 15899 3117
rect 15841 3077 15853 3111
rect 15887 3108 15899 3111
rect 18693 3111 18751 3117
rect 18693 3108 18705 3111
rect 15887 3080 18705 3108
rect 15887 3077 15899 3080
rect 15841 3071 15899 3077
rect 18693 3077 18705 3080
rect 18739 3108 18751 3111
rect 19886 3108 19892 3120
rect 18739 3080 19892 3108
rect 18739 3077 18751 3080
rect 18693 3071 18751 3077
rect 19886 3068 19892 3080
rect 19944 3068 19950 3120
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2924 3012 3065 3040
rect 2924 3000 2930 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3743 3012 3985 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8444 3012 8861 3040
rect 8444 3000 8450 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10192 3012 10885 3040
rect 10192 3000 10198 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 18506 3000 18512 3052
rect 18564 3000 18570 3052
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 7374 2972 7380 2984
rect 1903 2944 7380 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 1302 2864 1308 2916
rect 1360 2904 1366 2916
rect 1596 2904 1624 2935
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8076 2944 9137 2972
rect 8076 2932 8082 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 9824 2944 14289 2972
rect 9824 2932 9830 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2972 20407 2975
rect 22738 2972 22744 2984
rect 20395 2944 22744 2972
rect 20395 2941 20407 2944
rect 20349 2935 20407 2941
rect 22738 2932 22744 2944
rect 22796 2932 22802 2984
rect 4157 2907 4215 2913
rect 4157 2904 4169 2907
rect 1360 2876 4169 2904
rect 1360 2864 1366 2876
rect 4157 2873 4169 2876
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 2774 2836 2780 2848
rect 1452 2808 2780 2836
rect 1452 2796 1458 2808
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 4338 2796 4344 2848
rect 4396 2796 4402 2848
rect 11882 2796 11888 2848
rect 11940 2796 11946 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 15933 2839 15991 2845
rect 15933 2836 15945 2839
rect 12492 2808 15945 2836
rect 12492 2796 12498 2808
rect 15933 2805 15945 2808
rect 15979 2805 15991 2839
rect 15933 2799 15991 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 4338 2632 4344 2644
rect 1596 2604 4344 2632
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 1596 2505 1624 2604
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27522 2592 27528 2644
rect 27580 2632 27586 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27580 2604 28181 2632
rect 27580 2592 27586 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 29086 2592 29092 2644
rect 29144 2632 29150 2644
rect 30837 2635 30895 2641
rect 30837 2632 30849 2635
rect 29144 2604 30849 2632
rect 29144 2592 29150 2604
rect 30837 2601 30849 2604
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 33505 2635 33563 2641
rect 33505 2632 33517 2635
rect 32916 2604 33517 2632
rect 32916 2592 32922 2604
rect 33505 2601 33517 2604
rect 33551 2601 33563 2635
rect 33505 2595 33563 2601
rect 15010 2564 15016 2576
rect 1872 2536 15016 2564
rect 1872 2505 1900 2536
rect 15010 2524 15016 2536
rect 15068 2524 15074 2576
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1360 2468 1593 2496
rect 1360 2456 1366 2468
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2465 1915 2499
rect 2866 2496 2872 2508
rect 1857 2459 1915 2465
rect 2240 2468 2872 2496
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 2240 2428 2268 2468
rect 2866 2456 2872 2468
rect 2924 2496 2930 2508
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 2924 2468 3525 2496
rect 2924 2456 2930 2468
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 28718 2456 28724 2508
rect 28776 2496 28782 2508
rect 36357 2499 36415 2505
rect 36357 2496 36369 2499
rect 28776 2468 36369 2496
rect 28776 2456 28782 2468
rect 36357 2465 36369 2468
rect 36403 2465 36415 2499
rect 36357 2459 36415 2465
rect 1268 2400 2268 2428
rect 1268 2388 1274 2400
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2832 2400 3065 2428
rect 2832 2388 2838 2400
rect 3053 2397 3065 2400
rect 3099 2428 3111 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3099 2400 3801 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8294 2428 8300 2440
rect 7055 2400 8300 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 4356 2360 4384 2391
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 9766 2428 9772 2440
rect 9631 2400 9772 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12434 2428 12440 2440
rect 12391 2400 12440 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25731 2400 25973 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2428 33747 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33735 2400 33977 2428
rect 33735 2397 33747 2400
rect 33689 2391 33747 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 11882 2360 11888 2372
rect 3252 2332 4292 2360
rect 4356 2332 11888 2360
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 3252 2292 3280 2332
rect 2915 2264 3280 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 4264 2292 4292 2332
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 8018 2292 8024 2304
rect 4264 2264 8024 2292
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 1302 2048 1308 2100
rect 1360 2088 1366 2100
rect 3326 2088 3332 2100
rect 1360 2060 3332 2088
rect 1360 2048 1366 2060
rect 3326 2048 3332 2060
rect 3384 2048 3390 2100
<< via1 >>
rect 8852 26120 8904 26172
rect 30932 26120 30984 26172
rect 17868 26052 17920 26104
rect 33968 26052 34020 26104
rect 15016 25984 15068 26036
rect 35256 25984 35308 26036
rect 12440 25916 12492 25968
rect 36084 25916 36136 25968
rect 17408 25848 17460 25900
rect 40408 25848 40460 25900
rect 25044 25780 25096 25832
rect 39764 25780 39816 25832
rect 11796 25712 11848 25764
rect 36544 25712 36596 25764
rect 12256 25644 12308 25696
rect 38660 25644 38712 25696
rect 16672 25576 16724 25628
rect 36268 25576 36320 25628
rect 6276 25508 6328 25560
rect 35900 25508 35952 25560
rect 13544 25440 13596 25492
rect 33324 25440 33376 25492
rect 11060 25372 11112 25424
rect 34704 25372 34756 25424
rect 12072 25304 12124 25356
rect 34612 25304 34664 25356
rect 9864 25236 9916 25288
rect 32404 25236 32456 25288
rect 3884 25168 3936 25220
rect 9772 25168 9824 25220
rect 22560 25168 22612 25220
rect 32772 25168 32824 25220
rect 20628 25100 20680 25152
rect 32680 25100 32732 25152
rect 6644 25032 6696 25084
rect 22008 25032 22060 25084
rect 26148 25032 26200 25084
rect 39856 25032 39908 25084
rect 9128 24964 9180 25016
rect 17408 24964 17460 25016
rect 27160 24964 27212 25016
rect 40040 24964 40092 25016
rect 28908 24896 28960 24948
rect 35624 24896 35676 24948
rect 3148 24828 3200 24880
rect 4436 24828 4488 24880
rect 7104 24828 7156 24880
rect 15292 24828 15344 24880
rect 16672 24828 16724 24880
rect 29000 24828 29052 24880
rect 40132 24828 40184 24880
rect 14280 24760 14332 24812
rect 25504 24760 25556 24812
rect 26608 24760 26660 24812
rect 30104 24760 30156 24812
rect 35716 24760 35768 24812
rect 38384 24760 38436 24812
rect 4344 24692 4396 24744
rect 15016 24692 15068 24744
rect 15384 24692 15436 24744
rect 21180 24692 21232 24744
rect 27436 24692 27488 24744
rect 27528 24692 27580 24744
rect 29092 24692 29144 24744
rect 31208 24692 31260 24744
rect 37740 24692 37792 24744
rect 14924 24624 14976 24676
rect 24492 24624 24544 24676
rect 3792 24556 3844 24608
rect 21364 24556 21416 24608
rect 24400 24556 24452 24608
rect 29368 24624 29420 24676
rect 32220 24624 32272 24676
rect 36636 24624 36688 24676
rect 24860 24556 24912 24608
rect 27712 24556 27764 24608
rect 28080 24556 28132 24608
rect 29184 24556 29236 24608
rect 29276 24556 29328 24608
rect 36912 24556 36964 24608
rect 37004 24556 37056 24608
rect 39304 24556 39356 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 3976 24395 4028 24404
rect 3976 24361 3985 24395
rect 3985 24361 4019 24395
rect 4019 24361 4028 24395
rect 3976 24352 4028 24361
rect 4252 24352 4304 24404
rect 4344 24395 4396 24404
rect 4344 24361 4353 24395
rect 4353 24361 4387 24395
rect 4387 24361 4396 24395
rect 4344 24352 4396 24361
rect 24400 24352 24452 24404
rect 24492 24352 24544 24404
rect 25136 24352 25188 24404
rect 31576 24352 31628 24404
rect 32864 24352 32916 24404
rect 35072 24352 35124 24404
rect 39304 24395 39356 24404
rect 39304 24361 39313 24395
rect 39313 24361 39347 24395
rect 39347 24361 39356 24395
rect 39304 24352 39356 24361
rect 40040 24395 40092 24404
rect 40040 24361 40049 24395
rect 40049 24361 40083 24395
rect 40083 24361 40092 24395
rect 40040 24352 40092 24361
rect 44732 24395 44784 24404
rect 44732 24361 44741 24395
rect 44741 24361 44775 24395
rect 44775 24361 44784 24395
rect 44732 24352 44784 24361
rect 1584 24327 1636 24336
rect 1584 24293 1593 24327
rect 1593 24293 1627 24327
rect 1627 24293 1636 24327
rect 1584 24284 1636 24293
rect 2780 24284 2832 24336
rect 4712 24284 4764 24336
rect 9312 24284 9364 24336
rect 9404 24284 9456 24336
rect 3516 24216 3568 24268
rect 6828 24216 6880 24268
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 2136 24191 2188 24200
rect 2136 24157 2145 24191
rect 2145 24157 2179 24191
rect 2179 24157 2188 24191
rect 2136 24148 2188 24157
rect 756 24080 808 24132
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 9312 24191 9364 24200
rect 9312 24157 9321 24191
rect 9321 24157 9355 24191
rect 9355 24157 9364 24191
rect 9312 24148 9364 24157
rect 10048 24148 10100 24200
rect 3976 24080 4028 24132
rect 7472 24080 7524 24132
rect 8944 24080 8996 24132
rect 12624 24148 12676 24200
rect 14280 24327 14332 24336
rect 14280 24293 14289 24327
rect 14289 24293 14323 24327
rect 14323 24293 14332 24327
rect 14280 24284 14332 24293
rect 18880 24284 18932 24336
rect 23388 24284 23440 24336
rect 27620 24284 27672 24336
rect 29092 24284 29144 24336
rect 14372 24216 14424 24268
rect 14740 24216 14792 24268
rect 9496 24012 9548 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 13820 24080 13872 24132
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 14832 24148 14884 24200
rect 16028 24080 16080 24132
rect 16212 24080 16264 24132
rect 17132 24216 17184 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24216 21600 24268
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 25044 24216 25096 24268
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 26332 24259 26384 24268
rect 26332 24225 26341 24259
rect 26341 24225 26375 24259
rect 26375 24225 26384 24259
rect 26332 24216 26384 24225
rect 26976 24216 27028 24268
rect 28080 24216 28132 24268
rect 28356 24259 28408 24268
rect 28356 24225 28365 24259
rect 28365 24225 28399 24259
rect 28399 24225 28408 24259
rect 28356 24216 28408 24225
rect 29276 24216 29328 24268
rect 30564 24284 30616 24336
rect 31668 24216 31720 24268
rect 33048 24216 33100 24268
rect 25320 24148 25372 24200
rect 26148 24148 26200 24200
rect 26424 24148 26476 24200
rect 18420 24080 18472 24132
rect 19524 24080 19576 24132
rect 15384 24012 15436 24064
rect 15476 24012 15528 24064
rect 23664 24012 23716 24064
rect 24768 24012 24820 24064
rect 25688 24012 25740 24064
rect 26792 24080 26844 24132
rect 27804 24080 27856 24132
rect 28540 24080 28592 24132
rect 29092 24191 29144 24200
rect 29092 24157 29101 24191
rect 29101 24157 29135 24191
rect 29135 24157 29144 24191
rect 29092 24148 29144 24157
rect 29828 24148 29880 24200
rect 30104 24148 30156 24200
rect 31116 24148 31168 24200
rect 33876 24148 33928 24200
rect 34888 24191 34940 24200
rect 34888 24157 34897 24191
rect 34897 24157 34931 24191
rect 34931 24157 34940 24191
rect 34888 24148 34940 24157
rect 35808 24148 35860 24200
rect 33508 24080 33560 24132
rect 37372 24080 37424 24132
rect 38292 24148 38344 24200
rect 38660 24259 38712 24268
rect 38660 24225 38669 24259
rect 38669 24225 38703 24259
rect 38703 24225 38712 24259
rect 38660 24216 38712 24225
rect 43536 24284 43588 24336
rect 38936 24148 38988 24200
rect 39212 24191 39264 24200
rect 39212 24157 39221 24191
rect 39221 24157 39255 24191
rect 39255 24157 39264 24191
rect 39212 24148 39264 24157
rect 40316 24148 40368 24200
rect 41236 24191 41288 24200
rect 41236 24157 41245 24191
rect 41245 24157 41279 24191
rect 41279 24157 41288 24191
rect 41236 24148 41288 24157
rect 25964 24012 26016 24064
rect 26976 24055 27028 24064
rect 26976 24021 26985 24055
rect 26985 24021 27019 24055
rect 27019 24021 27028 24055
rect 26976 24012 27028 24021
rect 27252 24055 27304 24064
rect 27252 24021 27261 24055
rect 27261 24021 27295 24055
rect 27295 24021 27304 24055
rect 27252 24012 27304 24021
rect 27712 24055 27764 24064
rect 27712 24021 27721 24055
rect 27721 24021 27755 24055
rect 27755 24021 27764 24055
rect 27712 24012 27764 24021
rect 28080 24055 28132 24064
rect 28080 24021 28089 24055
rect 28089 24021 28123 24055
rect 28123 24021 28132 24055
rect 28080 24012 28132 24021
rect 28816 24012 28868 24064
rect 29000 24012 29052 24064
rect 32772 24012 32824 24064
rect 35808 24012 35860 24064
rect 35992 24012 36044 24064
rect 36728 24055 36780 24064
rect 36728 24021 36737 24055
rect 36737 24021 36771 24055
rect 36771 24021 36780 24055
rect 36728 24012 36780 24021
rect 37280 24012 37332 24064
rect 41512 24191 41564 24200
rect 41512 24157 41521 24191
rect 41521 24157 41555 24191
rect 41555 24157 41564 24191
rect 41512 24148 41564 24157
rect 41604 24148 41656 24200
rect 42616 24191 42668 24200
rect 42616 24157 42625 24191
rect 42625 24157 42659 24191
rect 42659 24157 42668 24191
rect 42616 24148 42668 24157
rect 44732 24148 44784 24200
rect 45560 24148 45612 24200
rect 46020 24148 46072 24200
rect 47308 24148 47360 24200
rect 47952 24148 48004 24200
rect 42432 24080 42484 24132
rect 42524 24080 42576 24132
rect 40776 24012 40828 24064
rect 43904 24055 43956 24064
rect 43904 24021 43913 24055
rect 43913 24021 43947 24055
rect 43947 24021 43956 24055
rect 43904 24012 43956 24021
rect 45284 24012 45336 24064
rect 47032 24012 47084 24064
rect 48596 24012 48648 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 9404 23808 9456 23860
rect 10140 23808 10192 23860
rect 15476 23808 15528 23860
rect 22284 23808 22336 23860
rect 22652 23808 22704 23860
rect 26976 23808 27028 23860
rect 2412 23740 2464 23792
rect 848 23604 900 23656
rect 4160 23672 4212 23724
rect 7656 23672 7708 23724
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 3700 23604 3752 23656
rect 4528 23604 4580 23656
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 7564 23604 7616 23656
rect 9956 23740 10008 23792
rect 12532 23740 12584 23792
rect 15752 23740 15804 23792
rect 19064 23740 19116 23792
rect 19248 23740 19300 23792
rect 20444 23740 20496 23792
rect 21364 23783 21416 23792
rect 21364 23749 21373 23783
rect 21373 23749 21407 23783
rect 21407 23749 21416 23783
rect 21364 23740 21416 23749
rect 23572 23740 23624 23792
rect 25136 23783 25188 23792
rect 25136 23749 25145 23783
rect 25145 23749 25179 23783
rect 25179 23749 25188 23783
rect 25136 23740 25188 23749
rect 26792 23740 26844 23792
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 10232 23604 10284 23656
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 13728 23672 13780 23724
rect 14372 23604 14424 23656
rect 14740 23672 14792 23724
rect 15016 23715 15068 23724
rect 15016 23681 15025 23715
rect 15025 23681 15059 23715
rect 15059 23681 15068 23715
rect 15016 23672 15068 23681
rect 16948 23672 17000 23724
rect 17408 23672 17460 23724
rect 21180 23715 21232 23724
rect 21180 23681 21189 23715
rect 21189 23681 21223 23715
rect 21223 23681 21232 23715
rect 21180 23672 21232 23681
rect 572 23468 624 23520
rect 2412 23468 2464 23520
rect 5540 23468 5592 23520
rect 6552 23468 6604 23520
rect 6644 23468 6696 23520
rect 9496 23468 9548 23520
rect 16304 23604 16356 23656
rect 20352 23604 20404 23656
rect 22652 23604 22704 23656
rect 22836 23604 22888 23656
rect 23296 23536 23348 23588
rect 25688 23604 25740 23656
rect 27436 23740 27488 23792
rect 27712 23740 27764 23792
rect 27896 23740 27948 23792
rect 28816 23808 28868 23860
rect 30196 23740 30248 23792
rect 30380 23740 30432 23792
rect 30748 23783 30800 23792
rect 30748 23749 30757 23783
rect 30757 23749 30791 23783
rect 30791 23749 30800 23783
rect 30748 23740 30800 23749
rect 32864 23808 32916 23860
rect 36544 23851 36596 23860
rect 36544 23817 36553 23851
rect 36553 23817 36587 23851
rect 36587 23817 36596 23851
rect 36544 23808 36596 23817
rect 36912 23851 36964 23860
rect 36912 23817 36921 23851
rect 36921 23817 36955 23851
rect 36955 23817 36964 23851
rect 36912 23808 36964 23817
rect 37464 23851 37516 23860
rect 37464 23817 37473 23851
rect 37473 23817 37507 23851
rect 37507 23817 37516 23851
rect 37464 23808 37516 23817
rect 38752 23808 38804 23860
rect 39212 23808 39264 23860
rect 42432 23851 42484 23860
rect 42432 23817 42441 23851
rect 42441 23817 42475 23851
rect 42475 23817 42484 23851
rect 42432 23808 42484 23817
rect 42616 23808 42668 23860
rect 43444 23808 43496 23860
rect 28724 23672 28776 23724
rect 30104 23672 30156 23724
rect 30932 23715 30984 23724
rect 30932 23681 30941 23715
rect 30941 23681 30975 23715
rect 30975 23681 30984 23715
rect 30932 23672 30984 23681
rect 31024 23672 31076 23724
rect 32220 23672 32272 23724
rect 34612 23715 34664 23724
rect 34612 23681 34621 23715
rect 34621 23681 34655 23715
rect 34655 23681 34664 23715
rect 34612 23672 34664 23681
rect 35716 23715 35768 23724
rect 26608 23579 26660 23588
rect 26608 23545 26617 23579
rect 26617 23545 26651 23579
rect 26651 23545 26660 23579
rect 26608 23536 26660 23545
rect 19708 23468 19760 23520
rect 19800 23468 19852 23520
rect 26424 23468 26476 23520
rect 29000 23604 29052 23656
rect 29368 23647 29420 23656
rect 29368 23613 29377 23647
rect 29377 23613 29411 23647
rect 29411 23613 29420 23647
rect 29368 23604 29420 23613
rect 30012 23604 30064 23656
rect 34336 23647 34388 23656
rect 34336 23613 34345 23647
rect 34345 23613 34379 23647
rect 34379 23613 34388 23647
rect 34336 23604 34388 23613
rect 34428 23604 34480 23656
rect 35716 23681 35742 23715
rect 35742 23681 35768 23715
rect 35716 23672 35768 23681
rect 35900 23715 35952 23724
rect 35900 23681 35909 23715
rect 35909 23681 35943 23715
rect 35943 23681 35952 23715
rect 35900 23672 35952 23681
rect 36452 23715 36504 23724
rect 36452 23681 36461 23715
rect 36461 23681 36495 23715
rect 36495 23681 36504 23715
rect 36452 23672 36504 23681
rect 36912 23672 36964 23724
rect 37740 23672 37792 23724
rect 40776 23740 40828 23792
rect 41236 23740 41288 23792
rect 45560 23808 45612 23860
rect 47308 23808 47360 23860
rect 39212 23672 39264 23724
rect 39948 23672 40000 23724
rect 40132 23672 40184 23724
rect 40408 23672 40460 23724
rect 35808 23604 35860 23656
rect 39580 23604 39632 23656
rect 44180 23672 44232 23724
rect 46664 23672 46716 23724
rect 48872 23715 48924 23724
rect 48872 23681 48881 23715
rect 48881 23681 48915 23715
rect 48915 23681 48924 23715
rect 48872 23672 48924 23681
rect 40960 23647 41012 23656
rect 40960 23613 40969 23647
rect 40969 23613 41003 23647
rect 41003 23613 41012 23647
rect 40960 23604 41012 23613
rect 41052 23604 41104 23656
rect 27528 23468 27580 23520
rect 27804 23468 27856 23520
rect 29276 23536 29328 23588
rect 31668 23536 31720 23588
rect 33876 23536 33928 23588
rect 31116 23468 31168 23520
rect 31392 23511 31444 23520
rect 31392 23477 31401 23511
rect 31401 23477 31435 23511
rect 31435 23477 31444 23511
rect 31392 23468 31444 23477
rect 31852 23511 31904 23520
rect 31852 23477 31861 23511
rect 31861 23477 31895 23511
rect 31895 23477 31904 23511
rect 31852 23468 31904 23477
rect 32220 23468 32272 23520
rect 33784 23511 33836 23520
rect 33784 23477 33793 23511
rect 33793 23477 33827 23511
rect 33827 23477 33836 23511
rect 33784 23468 33836 23477
rect 35624 23536 35676 23588
rect 38292 23536 38344 23588
rect 43444 23536 43496 23588
rect 40224 23468 40276 23520
rect 41052 23468 41104 23520
rect 43720 23511 43772 23520
rect 43720 23477 43729 23511
rect 43729 23477 43763 23511
rect 43763 23477 43772 23511
rect 43720 23468 43772 23477
rect 46940 23511 46992 23520
rect 46940 23477 46949 23511
rect 46949 23477 46983 23511
rect 46983 23477 46992 23511
rect 46940 23468 46992 23477
rect 48688 23511 48740 23520
rect 48688 23477 48697 23511
rect 48697 23477 48731 23511
rect 48731 23477 48740 23511
rect 48688 23468 48740 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 16212 23264 16264 23316
rect 18972 23264 19024 23316
rect 6828 23196 6880 23248
rect 9128 23239 9180 23248
rect 9128 23205 9137 23239
rect 9137 23205 9171 23239
rect 9171 23205 9180 23239
rect 9128 23196 9180 23205
rect 11152 23239 11204 23248
rect 11152 23205 11161 23239
rect 11161 23205 11195 23239
rect 11195 23205 11204 23239
rect 11152 23196 11204 23205
rect 23020 23264 23072 23316
rect 23112 23264 23164 23316
rect 21824 23239 21876 23248
rect 21824 23205 21833 23239
rect 21833 23205 21867 23239
rect 21867 23205 21876 23239
rect 21824 23196 21876 23205
rect 24676 23239 24728 23248
rect 24676 23205 24685 23239
rect 24685 23205 24719 23239
rect 24719 23205 24728 23239
rect 24676 23196 24728 23205
rect 5540 23128 5592 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 7012 23060 7064 23112
rect 7380 23060 7432 23112
rect 12532 23128 12584 23180
rect 9404 23103 9456 23112
rect 9404 23069 9413 23103
rect 9413 23069 9447 23103
rect 9447 23069 9456 23103
rect 9404 23060 9456 23069
rect 14556 23060 14608 23112
rect 17960 23128 18012 23180
rect 19708 23128 19760 23180
rect 20352 23128 20404 23180
rect 20444 23128 20496 23180
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 23296 23128 23348 23180
rect 23572 23128 23624 23180
rect 23756 23128 23808 23180
rect 30104 23264 30156 23316
rect 30196 23264 30248 23316
rect 28540 23196 28592 23248
rect 29092 23196 29144 23248
rect 32772 23264 32824 23316
rect 34980 23264 35032 23316
rect 37004 23264 37056 23316
rect 37096 23264 37148 23316
rect 34244 23196 34296 23248
rect 36452 23196 36504 23248
rect 26424 23171 26476 23180
rect 26424 23137 26433 23171
rect 26433 23137 26467 23171
rect 26467 23137 26476 23171
rect 26424 23128 26476 23137
rect 27252 23171 27304 23180
rect 27252 23137 27261 23171
rect 27261 23137 27295 23171
rect 27295 23137 27304 23171
rect 27252 23128 27304 23137
rect 28908 23128 28960 23180
rect 30012 23171 30064 23180
rect 30012 23137 30021 23171
rect 30021 23137 30055 23171
rect 30055 23137 30064 23171
rect 30012 23128 30064 23137
rect 32588 23128 32640 23180
rect 34796 23128 34848 23180
rect 23848 23060 23900 23112
rect 26056 23060 26108 23112
rect 26148 23060 26200 23112
rect 31760 23060 31812 23112
rect 31944 23103 31996 23112
rect 31944 23069 31953 23103
rect 31953 23069 31987 23103
rect 31987 23069 31996 23103
rect 31944 23060 31996 23069
rect 32036 23060 32088 23112
rect 32956 23060 33008 23112
rect 940 22924 992 22976
rect 5632 22992 5684 23044
rect 6460 22924 6512 22976
rect 9680 23035 9732 23044
rect 9680 23001 9689 23035
rect 9689 23001 9723 23035
rect 9723 23001 9732 23035
rect 9680 22992 9732 23001
rect 11428 22992 11480 23044
rect 11704 22992 11756 23044
rect 12072 22992 12124 23044
rect 13820 23035 13872 23044
rect 13820 23001 13829 23035
rect 13829 23001 13863 23035
rect 13863 23001 13872 23035
rect 13820 22992 13872 23001
rect 17316 22992 17368 23044
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 18420 22992 18472 23044
rect 20628 22992 20680 23044
rect 12624 22924 12676 22976
rect 12716 22924 12768 22976
rect 14556 22924 14608 22976
rect 16304 22924 16356 22976
rect 18328 22924 18380 22976
rect 22560 23035 22612 23044
rect 22560 23001 22569 23035
rect 22569 23001 22603 23035
rect 22603 23001 22612 23035
rect 22560 22992 22612 23001
rect 23572 22992 23624 23044
rect 26332 22992 26384 23044
rect 27436 22992 27488 23044
rect 29092 22992 29144 23044
rect 34336 23103 34388 23112
rect 34336 23069 34345 23103
rect 34345 23069 34379 23103
rect 34379 23069 34388 23103
rect 34336 23060 34388 23069
rect 35072 23103 35124 23112
rect 35072 23069 35081 23103
rect 35081 23069 35115 23103
rect 35115 23069 35124 23103
rect 35072 23060 35124 23069
rect 35532 23103 35584 23112
rect 35532 23069 35541 23103
rect 35541 23069 35575 23103
rect 35575 23069 35584 23103
rect 35532 23060 35584 23069
rect 35716 23128 35768 23180
rect 36912 23196 36964 23248
rect 37280 23196 37332 23248
rect 36728 23128 36780 23180
rect 40868 23196 40920 23248
rect 37004 23103 37056 23112
rect 37004 23069 37013 23103
rect 37013 23069 37047 23103
rect 37047 23069 37056 23103
rect 37004 23060 37056 23069
rect 37464 23060 37516 23112
rect 38476 23103 38528 23112
rect 38476 23069 38485 23103
rect 38485 23069 38519 23103
rect 38519 23069 38528 23103
rect 38476 23060 38528 23069
rect 38936 23103 38988 23112
rect 38936 23069 38945 23103
rect 38945 23069 38979 23103
rect 38979 23069 38988 23103
rect 38936 23060 38988 23069
rect 39764 23060 39816 23112
rect 40868 23103 40920 23112
rect 40868 23069 40877 23103
rect 40877 23069 40911 23103
rect 40911 23069 40920 23103
rect 40868 23060 40920 23069
rect 41144 23060 41196 23112
rect 24032 22967 24084 22976
rect 24032 22933 24041 22967
rect 24041 22933 24075 22967
rect 24075 22933 24084 22967
rect 24032 22924 24084 22933
rect 25136 22967 25188 22976
rect 25136 22933 25145 22967
rect 25145 22933 25179 22967
rect 25179 22933 25188 22967
rect 25136 22924 25188 22933
rect 25688 22924 25740 22976
rect 25964 22924 26016 22976
rect 26424 22924 26476 22976
rect 27712 22924 27764 22976
rect 30380 22924 30432 22976
rect 30656 22924 30708 22976
rect 31576 22924 31628 22976
rect 32956 22924 33008 22976
rect 34980 22992 35032 23044
rect 35164 22992 35216 23044
rect 37372 22992 37424 23044
rect 37556 23035 37608 23044
rect 37556 23001 37565 23035
rect 37565 23001 37599 23035
rect 37599 23001 37608 23035
rect 37556 22992 37608 23001
rect 38292 23035 38344 23044
rect 38292 23001 38301 23035
rect 38301 23001 38335 23035
rect 38335 23001 38344 23035
rect 38292 22992 38344 23001
rect 39580 22992 39632 23044
rect 33692 22967 33744 22976
rect 33692 22933 33701 22967
rect 33701 22933 33735 22967
rect 33735 22933 33744 22967
rect 33692 22924 33744 22933
rect 35900 22924 35952 22976
rect 37188 22924 37240 22976
rect 37648 22967 37700 22976
rect 37648 22933 37657 22967
rect 37657 22933 37691 22967
rect 37691 22933 37700 22967
rect 37648 22924 37700 22933
rect 39120 22967 39172 22976
rect 39120 22933 39129 22967
rect 39129 22933 39163 22967
rect 39163 22933 39172 22967
rect 39120 22924 39172 22933
rect 39856 22924 39908 22976
rect 41972 22967 42024 22976
rect 41972 22933 41981 22967
rect 41981 22933 42015 22967
rect 42015 22933 42024 22967
rect 41972 22924 42024 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 664 22720 716 22772
rect 5172 22652 5224 22704
rect 5264 22652 5316 22704
rect 7104 22695 7156 22704
rect 7104 22661 7113 22695
rect 7113 22661 7147 22695
rect 7147 22661 7156 22695
rect 7104 22652 7156 22661
rect 2872 22516 2924 22568
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 6920 22584 6972 22636
rect 9680 22720 9732 22772
rect 11060 22720 11112 22772
rect 12532 22720 12584 22772
rect 12624 22720 12676 22772
rect 14832 22720 14884 22772
rect 8576 22652 8628 22704
rect 5264 22448 5316 22500
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 10692 22695 10744 22704
rect 10692 22661 10701 22695
rect 10701 22661 10735 22695
rect 10735 22661 10744 22695
rect 10692 22652 10744 22661
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 11336 22584 11388 22636
rect 12716 22695 12768 22704
rect 12716 22661 12725 22695
rect 12725 22661 12759 22695
rect 12759 22661 12768 22695
rect 12716 22652 12768 22661
rect 13820 22584 13872 22636
rect 14924 22627 14976 22636
rect 14924 22593 14933 22627
rect 14933 22593 14967 22627
rect 14967 22593 14976 22627
rect 14924 22584 14976 22593
rect 10968 22516 11020 22568
rect 11152 22516 11204 22568
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 17224 22652 17276 22704
rect 18420 22652 18472 22704
rect 18880 22720 18932 22772
rect 19524 22652 19576 22704
rect 19984 22695 20036 22704
rect 19984 22661 19993 22695
rect 19993 22661 20027 22695
rect 20027 22661 20036 22695
rect 19984 22652 20036 22661
rect 20444 22652 20496 22704
rect 19708 22627 19760 22636
rect 19708 22593 19717 22627
rect 19717 22593 19751 22627
rect 19751 22593 19760 22627
rect 19708 22584 19760 22593
rect 23296 22652 23348 22704
rect 23480 22652 23532 22704
rect 23848 22652 23900 22704
rect 26332 22720 26384 22772
rect 27252 22720 27304 22772
rect 28908 22720 28960 22772
rect 31576 22763 31628 22772
rect 31576 22729 31585 22763
rect 31585 22729 31619 22763
rect 31619 22729 31628 22763
rect 31576 22720 31628 22729
rect 31668 22720 31720 22772
rect 33232 22720 33284 22772
rect 33876 22720 33928 22772
rect 5540 22380 5592 22432
rect 6460 22423 6512 22432
rect 6460 22389 6469 22423
rect 6469 22389 6503 22423
rect 6503 22389 6512 22423
rect 6460 22380 6512 22389
rect 11060 22380 11112 22432
rect 16764 22448 16816 22500
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 14188 22380 14240 22389
rect 14556 22423 14608 22432
rect 14556 22389 14565 22423
rect 14565 22389 14599 22423
rect 14599 22389 14608 22423
rect 14556 22380 14608 22389
rect 22744 22516 22796 22568
rect 23020 22516 23072 22568
rect 25228 22516 25280 22568
rect 30104 22652 30156 22704
rect 17132 22380 17184 22432
rect 18512 22380 18564 22432
rect 18972 22380 19024 22432
rect 23112 22448 23164 22500
rect 21456 22423 21508 22432
rect 21456 22389 21465 22423
rect 21465 22389 21499 22423
rect 21499 22389 21508 22423
rect 21456 22380 21508 22389
rect 23572 22380 23624 22432
rect 23756 22380 23808 22432
rect 25688 22448 25740 22500
rect 26056 22448 26108 22500
rect 27252 22516 27304 22568
rect 33692 22652 33744 22704
rect 34336 22720 34388 22772
rect 34428 22652 34480 22704
rect 36636 22652 36688 22704
rect 37372 22652 37424 22704
rect 40040 22720 40092 22772
rect 41144 22763 41196 22772
rect 41144 22729 41153 22763
rect 41153 22729 41187 22763
rect 41187 22729 41196 22763
rect 41144 22720 41196 22729
rect 39488 22652 39540 22704
rect 43904 22652 43956 22704
rect 31208 22584 31260 22636
rect 31852 22627 31904 22636
rect 31852 22593 31861 22627
rect 31861 22593 31895 22627
rect 31895 22593 31904 22627
rect 31852 22584 31904 22593
rect 32312 22627 32364 22636
rect 32312 22593 32321 22627
rect 32321 22593 32355 22627
rect 32355 22593 32364 22627
rect 32312 22584 32364 22593
rect 33876 22627 33928 22636
rect 33876 22593 33885 22627
rect 33885 22593 33919 22627
rect 33919 22593 33928 22627
rect 33876 22584 33928 22593
rect 34704 22584 34756 22636
rect 35624 22584 35676 22636
rect 36728 22584 36780 22636
rect 31024 22559 31076 22568
rect 31024 22525 31033 22559
rect 31033 22525 31067 22559
rect 31067 22525 31076 22559
rect 31024 22516 31076 22525
rect 31116 22559 31168 22568
rect 31116 22525 31125 22559
rect 31125 22525 31159 22559
rect 31159 22525 31168 22559
rect 31116 22516 31168 22525
rect 31576 22516 31628 22568
rect 33784 22516 33836 22568
rect 34336 22559 34388 22568
rect 34336 22525 34345 22559
rect 34345 22525 34379 22559
rect 34379 22525 34388 22559
rect 34336 22516 34388 22525
rect 35992 22516 36044 22568
rect 27620 22448 27672 22500
rect 30380 22448 30432 22500
rect 30840 22448 30892 22500
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 25780 22380 25832 22432
rect 26516 22380 26568 22432
rect 26608 22423 26660 22432
rect 26608 22389 26617 22423
rect 26617 22389 26651 22423
rect 26651 22389 26660 22423
rect 26608 22380 26660 22389
rect 27804 22423 27856 22432
rect 27804 22389 27813 22423
rect 27813 22389 27847 22423
rect 27847 22389 27856 22423
rect 27804 22380 27856 22389
rect 29184 22380 29236 22432
rect 30104 22423 30156 22432
rect 30104 22389 30113 22423
rect 30113 22389 30147 22423
rect 30147 22389 30156 22423
rect 30104 22380 30156 22389
rect 30196 22380 30248 22432
rect 31760 22380 31812 22432
rect 32036 22380 32088 22432
rect 33232 22380 33284 22432
rect 33600 22448 33652 22500
rect 37832 22516 37884 22568
rect 48688 22516 48740 22568
rect 35900 22380 35952 22432
rect 36084 22380 36136 22432
rect 36912 22423 36964 22432
rect 36912 22389 36921 22423
rect 36921 22389 36955 22423
rect 36955 22389 36964 22423
rect 36912 22380 36964 22389
rect 38384 22380 38436 22432
rect 40868 22448 40920 22500
rect 39764 22380 39816 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 4068 22176 4120 22228
rect 6644 22176 6696 22228
rect 9772 22176 9824 22228
rect 11152 22176 11204 22228
rect 11336 22176 11388 22228
rect 16304 22176 16356 22228
rect 17868 22176 17920 22228
rect 19340 22176 19392 22228
rect 20444 22176 20496 22228
rect 21456 22176 21508 22228
rect 25136 22176 25188 22228
rect 27804 22176 27856 22228
rect 28908 22176 28960 22228
rect 3792 22108 3844 22160
rect 5540 22108 5592 22160
rect 1308 22040 1360 22092
rect 3700 22040 3752 22092
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 6920 22108 6972 22160
rect 4160 21904 4212 21956
rect 7564 22040 7616 22092
rect 7840 22040 7892 22092
rect 10692 22108 10744 22160
rect 10876 22108 10928 22160
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 9956 22083 10008 22092
rect 9956 22049 9965 22083
rect 9965 22049 9999 22083
rect 9999 22049 10008 22083
rect 9956 22040 10008 22049
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 5632 21947 5684 21956
rect 5632 21913 5641 21947
rect 5641 21913 5675 21947
rect 5675 21913 5684 21947
rect 5632 21904 5684 21913
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 4344 21836 4396 21888
rect 5908 21879 5960 21888
rect 5908 21845 5917 21879
rect 5917 21845 5951 21879
rect 5951 21845 5960 21879
rect 5908 21836 5960 21845
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 10508 21972 10560 22024
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 10876 21972 10928 22024
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 13912 22108 13964 22160
rect 14556 22108 14608 22160
rect 15108 22108 15160 22160
rect 20628 22108 20680 22160
rect 21824 22108 21876 22160
rect 23296 22151 23348 22160
rect 23296 22117 23305 22151
rect 23305 22117 23339 22151
rect 23339 22117 23348 22151
rect 23296 22108 23348 22117
rect 13084 21972 13136 22024
rect 19432 22040 19484 22092
rect 19708 22040 19760 22092
rect 20536 22040 20588 22092
rect 25780 22108 25832 22160
rect 28356 22108 28408 22160
rect 31944 22176 31996 22228
rect 32496 22176 32548 22228
rect 36268 22176 36320 22228
rect 38292 22176 38344 22228
rect 30564 22108 30616 22160
rect 31116 22108 31168 22160
rect 34428 22108 34480 22160
rect 39488 22176 39540 22228
rect 7748 21904 7800 21956
rect 8852 21904 8904 21956
rect 8300 21836 8352 21888
rect 9220 21836 9272 21888
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 10600 21836 10652 21888
rect 11060 21904 11112 21956
rect 15568 21972 15620 22024
rect 18788 21972 18840 22024
rect 22652 21972 22704 22024
rect 23664 22015 23716 22024
rect 23664 21981 23673 22015
rect 23673 21981 23707 22015
rect 23707 21981 23716 22015
rect 23664 21972 23716 21981
rect 24860 22040 24912 22092
rect 25136 22040 25188 22092
rect 24308 21972 24360 22024
rect 27804 21972 27856 22024
rect 14096 21904 14148 21956
rect 14280 21836 14332 21888
rect 14648 21879 14700 21888
rect 14648 21845 14657 21879
rect 14657 21845 14691 21879
rect 14691 21845 14700 21879
rect 14648 21836 14700 21845
rect 14924 21836 14976 21888
rect 15108 21836 15160 21888
rect 16120 21836 16172 21888
rect 17868 21904 17920 21956
rect 19524 21947 19576 21956
rect 19524 21913 19533 21947
rect 19533 21913 19567 21947
rect 19567 21913 19576 21947
rect 19524 21904 19576 21913
rect 18880 21879 18932 21888
rect 18880 21845 18889 21879
rect 18889 21845 18923 21879
rect 18923 21845 18932 21879
rect 18880 21836 18932 21845
rect 19248 21836 19300 21888
rect 19340 21836 19392 21888
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 20076 21836 20128 21888
rect 24492 21836 24544 21888
rect 25504 21904 25556 21956
rect 25596 21904 25648 21956
rect 26056 21904 26108 21956
rect 26516 21904 26568 21956
rect 27344 21904 27396 21956
rect 29184 21904 29236 21956
rect 29368 22040 29420 22092
rect 30288 22040 30340 22092
rect 30656 22083 30708 22092
rect 30656 22049 30665 22083
rect 30665 22049 30699 22083
rect 30699 22049 30708 22083
rect 30656 22040 30708 22049
rect 31024 22040 31076 22092
rect 30104 21972 30156 22024
rect 32772 22040 32824 22092
rect 35256 22040 35308 22092
rect 36268 22040 36320 22092
rect 31944 21904 31996 21956
rect 33876 21904 33928 21956
rect 24952 21879 25004 21888
rect 24952 21845 24961 21879
rect 24961 21845 24995 21879
rect 24995 21845 25004 21879
rect 24952 21836 25004 21845
rect 26240 21836 26292 21888
rect 29092 21879 29144 21888
rect 29092 21845 29101 21879
rect 29101 21845 29135 21879
rect 29135 21845 29144 21879
rect 29092 21836 29144 21845
rect 29368 21836 29420 21888
rect 30012 21879 30064 21888
rect 30012 21845 30021 21879
rect 30021 21845 30055 21879
rect 30055 21845 30064 21879
rect 30012 21836 30064 21845
rect 30288 21836 30340 21888
rect 30472 21836 30524 21888
rect 32128 21836 32180 21888
rect 34612 21904 34664 21956
rect 35716 21947 35768 21956
rect 35716 21913 35725 21947
rect 35725 21913 35759 21947
rect 35759 21913 35768 21947
rect 35716 21904 35768 21913
rect 35900 21947 35952 21956
rect 35900 21913 35909 21947
rect 35909 21913 35943 21947
rect 35943 21913 35952 21947
rect 35900 21904 35952 21913
rect 37096 22015 37148 22024
rect 37096 21981 37105 22015
rect 37105 21981 37139 22015
rect 37139 21981 37148 22015
rect 37096 21972 37148 21981
rect 37740 22015 37792 22024
rect 37740 21981 37749 22015
rect 37749 21981 37783 22015
rect 37783 21981 37792 22015
rect 37740 21972 37792 21981
rect 37924 21972 37976 22024
rect 38292 21972 38344 22024
rect 39856 22040 39908 22092
rect 36268 21836 36320 21888
rect 37096 21836 37148 21888
rect 37188 21836 37240 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 4160 21632 4212 21684
rect 6920 21632 6972 21684
rect 8484 21632 8536 21684
rect 3240 21564 3292 21616
rect 3700 21564 3752 21616
rect 2320 21496 2372 21548
rect 3332 21428 3384 21480
rect 3608 21428 3660 21480
rect 6092 21428 6144 21480
rect 1124 21360 1176 21412
rect 3240 21292 3292 21344
rect 3424 21292 3476 21344
rect 4988 21292 5040 21344
rect 5448 21292 5500 21344
rect 7196 21471 7248 21480
rect 7196 21437 7205 21471
rect 7205 21437 7239 21471
rect 7239 21437 7248 21471
rect 7196 21428 7248 21437
rect 7104 21360 7156 21412
rect 7564 21360 7616 21412
rect 8116 21607 8168 21616
rect 8116 21573 8125 21607
rect 8125 21573 8159 21607
rect 8159 21573 8168 21607
rect 8116 21564 8168 21573
rect 9128 21564 9180 21616
rect 10876 21632 10928 21684
rect 10968 21632 11020 21684
rect 12440 21632 12492 21684
rect 11796 21564 11848 21616
rect 12532 21564 12584 21616
rect 14280 21632 14332 21684
rect 9772 21496 9824 21548
rect 11612 21496 11664 21548
rect 7840 21471 7892 21480
rect 7840 21437 7849 21471
rect 7849 21437 7883 21471
rect 7883 21437 7892 21471
rect 7840 21428 7892 21437
rect 10324 21428 10376 21480
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 12164 21428 12216 21480
rect 13728 21564 13780 21616
rect 14924 21564 14976 21616
rect 18788 21564 18840 21616
rect 19340 21564 19392 21616
rect 23204 21564 23256 21616
rect 23572 21564 23624 21616
rect 23940 21564 23992 21616
rect 25044 21632 25096 21684
rect 26148 21632 26200 21684
rect 28632 21632 28684 21684
rect 25320 21564 25372 21616
rect 30012 21632 30064 21684
rect 30656 21675 30708 21684
rect 30656 21641 30665 21675
rect 30665 21641 30699 21675
rect 30699 21641 30708 21675
rect 30656 21632 30708 21641
rect 31024 21675 31076 21684
rect 31024 21641 31033 21675
rect 31033 21641 31067 21675
rect 31067 21641 31076 21675
rect 31024 21632 31076 21641
rect 33232 21632 33284 21684
rect 33416 21675 33468 21684
rect 33416 21641 33425 21675
rect 33425 21641 33459 21675
rect 33459 21641 33468 21675
rect 33416 21632 33468 21641
rect 34704 21675 34756 21684
rect 34704 21641 34713 21675
rect 34713 21641 34747 21675
rect 34747 21641 34756 21675
rect 34704 21632 34756 21641
rect 36176 21632 36228 21684
rect 36820 21632 36872 21684
rect 37832 21632 37884 21684
rect 29368 21564 29420 21616
rect 30748 21564 30800 21616
rect 34336 21564 34388 21616
rect 14556 21496 14608 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 17776 21496 17828 21548
rect 18512 21496 18564 21548
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 20904 21496 20956 21548
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 25044 21496 25096 21548
rect 27252 21496 27304 21548
rect 27528 21496 27580 21548
rect 27712 21496 27764 21548
rect 28356 21496 28408 21548
rect 30288 21496 30340 21548
rect 32220 21496 32272 21548
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32772 21496 32824 21548
rect 12808 21428 12860 21480
rect 13544 21428 13596 21480
rect 14004 21428 14056 21480
rect 16028 21471 16080 21480
rect 16028 21437 16037 21471
rect 16037 21437 16071 21471
rect 16071 21437 16080 21471
rect 16028 21428 16080 21437
rect 6920 21292 6972 21344
rect 10784 21360 10836 21412
rect 11520 21360 11572 21412
rect 12716 21360 12768 21412
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 17132 21428 17184 21480
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 11428 21292 11480 21344
rect 13544 21292 13596 21344
rect 17684 21360 17736 21412
rect 17776 21360 17828 21412
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 27344 21428 27396 21480
rect 27804 21471 27856 21480
rect 27804 21437 27813 21471
rect 27813 21437 27847 21471
rect 27847 21437 27856 21471
rect 27804 21428 27856 21437
rect 15568 21335 15620 21344
rect 15568 21301 15577 21335
rect 15577 21301 15611 21335
rect 15611 21301 15620 21335
rect 15568 21292 15620 21301
rect 17224 21292 17276 21344
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 17500 21292 17552 21344
rect 22284 21360 22336 21412
rect 22376 21360 22428 21412
rect 20720 21292 20772 21344
rect 21456 21335 21508 21344
rect 21456 21301 21465 21335
rect 21465 21301 21499 21335
rect 21499 21301 21508 21335
rect 21456 21292 21508 21301
rect 21548 21292 21600 21344
rect 23388 21292 23440 21344
rect 26700 21403 26752 21412
rect 26700 21369 26709 21403
rect 26709 21369 26743 21403
rect 26743 21369 26752 21403
rect 30472 21428 30524 21480
rect 26700 21360 26752 21369
rect 25964 21292 26016 21344
rect 26976 21292 27028 21344
rect 30840 21360 30892 21412
rect 28908 21292 28960 21344
rect 29092 21292 29144 21344
rect 31024 21292 31076 21344
rect 34888 21496 34940 21548
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 35532 21564 35584 21616
rect 38292 21607 38344 21616
rect 38292 21573 38301 21607
rect 38301 21573 38335 21607
rect 38335 21573 38344 21607
rect 38292 21564 38344 21573
rect 36268 21496 36320 21548
rect 36360 21496 36412 21548
rect 47584 21496 47636 21548
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 32036 21360 32088 21412
rect 32220 21360 32272 21412
rect 32128 21292 32180 21344
rect 33232 21360 33284 21412
rect 36728 21360 36780 21412
rect 34612 21292 34664 21344
rect 36912 21292 36964 21344
rect 37832 21292 37884 21344
rect 47584 21335 47636 21344
rect 47584 21301 47593 21335
rect 47593 21301 47627 21335
rect 47627 21301 47636 21335
rect 47584 21292 47636 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 3792 21088 3844 21140
rect 3976 21088 4028 21140
rect 5816 21131 5868 21140
rect 5816 21097 5825 21131
rect 5825 21097 5859 21131
rect 5859 21097 5868 21131
rect 5816 21088 5868 21097
rect 5908 21088 5960 21140
rect 6000 21020 6052 21072
rect 8024 21131 8076 21140
rect 8024 21097 8033 21131
rect 8033 21097 8067 21131
rect 8067 21097 8076 21131
rect 8024 21088 8076 21097
rect 16028 21088 16080 21140
rect 16120 21088 16172 21140
rect 13544 21020 13596 21072
rect 13912 21020 13964 21072
rect 3516 20952 3568 21004
rect 7840 20952 7892 21004
rect 7932 20952 7984 21004
rect 11520 20952 11572 21004
rect 11888 20952 11940 21004
rect 2872 20816 2924 20868
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 9496 20884 9548 20936
rect 480 20748 532 20800
rect 3608 20791 3660 20800
rect 3608 20757 3617 20791
rect 3617 20757 3651 20791
rect 3651 20757 3660 20791
rect 3608 20748 3660 20757
rect 4160 20816 4212 20868
rect 5908 20791 5960 20800
rect 5908 20757 5917 20791
rect 5917 20757 5951 20791
rect 5951 20757 5960 20791
rect 5908 20748 5960 20757
rect 6552 20859 6604 20868
rect 6552 20825 6561 20859
rect 6561 20825 6595 20859
rect 6595 20825 6604 20859
rect 6552 20816 6604 20825
rect 7564 20816 7616 20868
rect 9680 20816 9732 20868
rect 12348 20884 12400 20936
rect 13452 20952 13504 21004
rect 14096 20952 14148 21004
rect 12716 20884 12768 20936
rect 14280 20995 14332 21004
rect 14280 20961 14289 20995
rect 14289 20961 14323 20995
rect 14323 20961 14332 20995
rect 14280 20952 14332 20961
rect 14924 20952 14976 21004
rect 15016 20952 15068 21004
rect 15660 20952 15712 21004
rect 17408 21020 17460 21072
rect 16488 20995 16540 21004
rect 16488 20961 16497 20995
rect 16497 20961 16531 20995
rect 16531 20961 16540 20995
rect 16488 20952 16540 20961
rect 17040 20952 17092 21004
rect 21824 21088 21876 21140
rect 22284 21088 22336 21140
rect 20720 21020 20772 21072
rect 19340 20952 19392 21004
rect 19432 20995 19484 21004
rect 19432 20961 19441 20995
rect 19441 20961 19475 20995
rect 19475 20961 19484 20995
rect 19432 20952 19484 20961
rect 20168 20952 20220 21004
rect 22468 20952 22520 21004
rect 23664 20995 23716 21004
rect 23664 20961 23673 20995
rect 23673 20961 23707 20995
rect 23707 20961 23716 20995
rect 23664 20952 23716 20961
rect 25964 21020 26016 21072
rect 27528 21088 27580 21140
rect 28908 21088 28960 21140
rect 31760 21088 31812 21140
rect 32036 21088 32088 21140
rect 33968 21088 34020 21140
rect 37372 21131 37424 21140
rect 37372 21097 37381 21131
rect 37381 21097 37415 21131
rect 37415 21097 37424 21131
rect 37372 21088 37424 21097
rect 30656 21020 30708 21072
rect 32404 21020 32456 21072
rect 14832 20884 14884 20936
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 18512 20884 18564 20936
rect 19248 20884 19300 20936
rect 24308 20884 24360 20936
rect 26700 20952 26752 21004
rect 26976 20952 27028 21004
rect 28448 20884 28500 20936
rect 28540 20884 28592 20936
rect 29092 20884 29144 20936
rect 29368 20884 29420 20936
rect 30196 20884 30248 20936
rect 30840 20927 30892 20936
rect 30840 20893 30849 20927
rect 30849 20893 30883 20927
rect 30883 20893 30892 20927
rect 30840 20884 30892 20893
rect 8392 20748 8444 20800
rect 8576 20748 8628 20800
rect 11152 20791 11204 20800
rect 11152 20757 11161 20791
rect 11161 20757 11195 20791
rect 11195 20757 11204 20791
rect 11152 20748 11204 20757
rect 17224 20816 17276 20868
rect 12256 20748 12308 20800
rect 12348 20748 12400 20800
rect 13912 20748 13964 20800
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 16396 20748 16448 20800
rect 18788 20791 18840 20800
rect 18788 20757 18797 20791
rect 18797 20757 18831 20791
rect 18831 20757 18840 20791
rect 18788 20748 18840 20757
rect 19616 20816 19668 20868
rect 19432 20748 19484 20800
rect 19984 20816 20036 20868
rect 21640 20859 21692 20868
rect 21640 20825 21649 20859
rect 21649 20825 21683 20859
rect 21683 20825 21692 20859
rect 21640 20816 21692 20825
rect 21824 20816 21876 20868
rect 23756 20816 23808 20868
rect 23940 20816 23992 20868
rect 24860 20816 24912 20868
rect 20352 20748 20404 20800
rect 21088 20748 21140 20800
rect 23572 20748 23624 20800
rect 24308 20748 24360 20800
rect 24584 20748 24636 20800
rect 25596 20748 25648 20800
rect 26240 20859 26292 20868
rect 26240 20825 26249 20859
rect 26249 20825 26283 20859
rect 26283 20825 26292 20859
rect 26240 20816 26292 20825
rect 26516 20816 26568 20868
rect 32864 20995 32916 21004
rect 32864 20961 32873 20995
rect 32873 20961 32907 20995
rect 32907 20961 32916 20995
rect 32864 20952 32916 20961
rect 33324 20952 33376 21004
rect 34336 20927 34388 20936
rect 34336 20893 34345 20927
rect 34345 20893 34379 20927
rect 34379 20893 34388 20927
rect 34336 20884 34388 20893
rect 36636 20884 36688 20936
rect 46848 20884 46900 20936
rect 35256 20816 35308 20868
rect 35440 20816 35492 20868
rect 36452 20859 36504 20868
rect 36452 20825 36461 20859
rect 36461 20825 36495 20859
rect 36495 20825 36504 20859
rect 36452 20816 36504 20825
rect 28816 20791 28868 20800
rect 28816 20757 28825 20791
rect 28825 20757 28859 20791
rect 28859 20757 28868 20791
rect 28816 20748 28868 20757
rect 29184 20748 29236 20800
rect 31484 20791 31536 20800
rect 31484 20757 31493 20791
rect 31493 20757 31527 20791
rect 31527 20757 31536 20791
rect 31484 20748 31536 20757
rect 35072 20791 35124 20800
rect 35072 20757 35081 20791
rect 35081 20757 35115 20791
rect 35115 20757 35124 20791
rect 35072 20748 35124 20757
rect 36544 20791 36596 20800
rect 36544 20757 36553 20791
rect 36553 20757 36587 20791
rect 36587 20757 36596 20791
rect 36544 20748 36596 20757
rect 37096 20791 37148 20800
rect 37096 20757 37105 20791
rect 37105 20757 37139 20791
rect 37139 20757 37148 20791
rect 37096 20748 37148 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 1032 20544 1084 20596
rect 5264 20544 5316 20596
rect 6460 20544 6512 20596
rect 1952 20408 2004 20460
rect 6184 20476 6236 20528
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 5632 20408 5684 20460
rect 6368 20408 6420 20460
rect 2412 20272 2464 20324
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5540 20340 5592 20392
rect 5908 20340 5960 20392
rect 6644 20340 6696 20392
rect 3700 20272 3752 20324
rect 11980 20587 12032 20596
rect 11980 20553 11989 20587
rect 11989 20553 12023 20587
rect 12023 20553 12032 20587
rect 11980 20544 12032 20553
rect 15568 20544 15620 20596
rect 16672 20587 16724 20596
rect 16672 20553 16681 20587
rect 16681 20553 16715 20587
rect 16715 20553 16724 20587
rect 16672 20544 16724 20553
rect 16948 20544 17000 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 7564 20340 7616 20392
rect 9128 20476 9180 20528
rect 11244 20476 11296 20528
rect 11704 20476 11756 20528
rect 12808 20476 12860 20528
rect 13636 20476 13688 20528
rect 14004 20519 14056 20528
rect 14004 20485 14013 20519
rect 14013 20485 14047 20519
rect 14047 20485 14056 20519
rect 14004 20476 14056 20485
rect 14280 20476 14332 20528
rect 14556 20476 14608 20528
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 17776 20476 17828 20528
rect 20720 20476 20772 20528
rect 10692 20408 10744 20460
rect 7288 20272 7340 20324
rect 7840 20272 7892 20324
rect 8852 20383 8904 20392
rect 8852 20349 8861 20383
rect 8861 20349 8895 20383
rect 8895 20349 8904 20383
rect 8852 20340 8904 20349
rect 9496 20340 9548 20392
rect 10876 20340 10928 20392
rect 13544 20408 13596 20460
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 17868 20408 17920 20460
rect 18788 20408 18840 20460
rect 13360 20340 13412 20392
rect 14096 20340 14148 20392
rect 5724 20204 5776 20256
rect 5816 20204 5868 20256
rect 8208 20204 8260 20256
rect 9956 20272 10008 20324
rect 9404 20204 9456 20256
rect 9864 20204 9916 20256
rect 11060 20204 11112 20256
rect 11428 20204 11480 20256
rect 12348 20204 12400 20256
rect 12716 20204 12768 20256
rect 15200 20204 15252 20256
rect 17684 20340 17736 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 19616 20408 19668 20460
rect 23572 20587 23624 20596
rect 23572 20553 23581 20587
rect 23581 20553 23615 20587
rect 23615 20553 23624 20587
rect 23572 20544 23624 20553
rect 23848 20544 23900 20596
rect 27436 20544 27488 20596
rect 23388 20476 23440 20528
rect 23388 20340 23440 20392
rect 19708 20272 19760 20324
rect 20996 20272 21048 20324
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 17132 20204 17184 20256
rect 18236 20204 18288 20256
rect 18420 20204 18472 20256
rect 18696 20204 18748 20256
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 23756 20383 23808 20392
rect 23756 20349 23765 20383
rect 23765 20349 23799 20383
rect 23799 20349 23808 20383
rect 23756 20340 23808 20349
rect 24492 20476 24544 20528
rect 24860 20476 24912 20528
rect 26516 20476 26568 20528
rect 26884 20476 26936 20528
rect 26976 20476 27028 20528
rect 27528 20451 27580 20460
rect 24308 20383 24360 20392
rect 24308 20349 24317 20383
rect 24317 20349 24351 20383
rect 24351 20349 24360 20383
rect 24308 20340 24360 20349
rect 25320 20340 25372 20392
rect 27528 20417 27537 20451
rect 27537 20417 27571 20451
rect 27571 20417 27580 20451
rect 27528 20408 27580 20417
rect 27160 20340 27212 20392
rect 31484 20544 31536 20596
rect 31760 20587 31812 20596
rect 31760 20553 31769 20587
rect 31769 20553 31803 20587
rect 31803 20553 31812 20587
rect 31760 20544 31812 20553
rect 31852 20587 31904 20596
rect 31852 20553 31861 20587
rect 31861 20553 31895 20587
rect 31895 20553 31904 20587
rect 31852 20544 31904 20553
rect 32864 20544 32916 20596
rect 34980 20544 35032 20596
rect 29368 20476 29420 20528
rect 27988 20408 28040 20460
rect 28356 20408 28408 20460
rect 26976 20272 27028 20324
rect 30196 20383 30248 20392
rect 30196 20349 30205 20383
rect 30205 20349 30239 20383
rect 30239 20349 30248 20383
rect 30196 20340 30248 20349
rect 28080 20272 28132 20324
rect 24768 20204 24820 20256
rect 26240 20204 26292 20256
rect 27528 20204 27580 20256
rect 30380 20272 30432 20324
rect 31208 20383 31260 20392
rect 31208 20349 31217 20383
rect 31217 20349 31251 20383
rect 31251 20349 31260 20383
rect 31208 20340 31260 20349
rect 31852 20272 31904 20324
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 32680 20476 32732 20528
rect 35532 20544 35584 20596
rect 39580 20476 39632 20528
rect 33692 20451 33744 20460
rect 33692 20417 33701 20451
rect 33701 20417 33735 20451
rect 33735 20417 33744 20451
rect 33692 20408 33744 20417
rect 40960 20408 41012 20460
rect 34980 20272 35032 20324
rect 35164 20272 35216 20324
rect 35624 20340 35676 20392
rect 35348 20272 35400 20324
rect 35716 20272 35768 20324
rect 29920 20204 29972 20256
rect 32036 20204 32088 20256
rect 33784 20247 33836 20256
rect 33784 20213 33793 20247
rect 33793 20213 33827 20247
rect 33827 20213 33836 20247
rect 33784 20204 33836 20213
rect 34520 20247 34572 20256
rect 34520 20213 34529 20247
rect 34529 20213 34563 20247
rect 34563 20213 34572 20247
rect 34520 20204 34572 20213
rect 35256 20247 35308 20256
rect 35256 20213 35265 20247
rect 35265 20213 35299 20247
rect 35299 20213 35308 20247
rect 35256 20204 35308 20213
rect 35440 20247 35492 20256
rect 35440 20213 35449 20247
rect 35449 20213 35483 20247
rect 35483 20213 35492 20247
rect 35440 20204 35492 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3608 20043 3660 20052
rect 3608 20009 3617 20043
rect 3617 20009 3651 20043
rect 3651 20009 3660 20043
rect 3608 20000 3660 20009
rect 4160 20043 4212 20052
rect 4160 20009 4169 20043
rect 4169 20009 4203 20043
rect 4203 20009 4212 20043
rect 4160 20000 4212 20009
rect 6920 20000 6972 20052
rect 8208 20000 8260 20052
rect 11612 20000 11664 20052
rect 7840 19932 7892 19984
rect 9496 19932 9548 19984
rect 11336 19932 11388 19984
rect 14096 20000 14148 20052
rect 14556 20000 14608 20052
rect 15016 20000 15068 20052
rect 15568 20000 15620 20052
rect 7380 19864 7432 19916
rect 7472 19864 7524 19916
rect 2504 19796 2556 19848
rect 2872 19728 2924 19780
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 9956 19864 10008 19916
rect 13728 19932 13780 19984
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 17132 19932 17184 19984
rect 9404 19839 9456 19848
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 11612 19796 11664 19848
rect 4528 19728 4580 19780
rect 5632 19728 5684 19780
rect 8300 19728 8352 19780
rect 5816 19660 5868 19712
rect 6000 19660 6052 19712
rect 6736 19660 6788 19712
rect 10048 19728 10100 19780
rect 11060 19728 11112 19780
rect 12348 19771 12400 19780
rect 12348 19737 12357 19771
rect 12357 19737 12391 19771
rect 12391 19737 12400 19771
rect 12348 19728 12400 19737
rect 12808 19728 12860 19780
rect 14096 19796 14148 19848
rect 17132 19796 17184 19848
rect 17960 19864 18012 19916
rect 18236 19932 18288 19984
rect 19432 19932 19484 19984
rect 20628 20000 20680 20052
rect 21916 20043 21968 20052
rect 21916 20009 21925 20043
rect 21925 20009 21959 20043
rect 21959 20009 21968 20043
rect 21916 20000 21968 20009
rect 25964 20000 26016 20052
rect 27804 20000 27856 20052
rect 27896 20000 27948 20052
rect 28816 19932 28868 19984
rect 28908 19932 28960 19984
rect 31300 19932 31352 19984
rect 19616 19864 19668 19916
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 22652 19864 22704 19916
rect 25044 19864 25096 19916
rect 25320 19907 25372 19916
rect 25320 19873 25329 19907
rect 25329 19873 25363 19907
rect 25363 19873 25372 19907
rect 25320 19864 25372 19873
rect 25780 19864 25832 19916
rect 27620 19864 27672 19916
rect 27712 19864 27764 19916
rect 20076 19796 20128 19848
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 22744 19796 22796 19848
rect 15016 19728 15068 19780
rect 11336 19660 11388 19712
rect 12256 19660 12308 19712
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 13544 19660 13596 19712
rect 14004 19660 14056 19712
rect 16672 19728 16724 19780
rect 18328 19728 18380 19780
rect 16488 19660 16540 19712
rect 19892 19728 19944 19780
rect 20352 19728 20404 19780
rect 20720 19728 20772 19780
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 19800 19660 19852 19712
rect 21088 19660 21140 19712
rect 22928 19660 22980 19712
rect 23664 19660 23716 19712
rect 24308 19660 24360 19712
rect 25228 19728 25280 19780
rect 27988 19796 28040 19848
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 29092 19864 29144 19916
rect 29276 19864 29328 19916
rect 30380 19796 30432 19848
rect 34336 20000 34388 20052
rect 31484 19864 31536 19916
rect 31668 19864 31720 19916
rect 33600 19864 33652 19916
rect 26148 19728 26200 19780
rect 26884 19728 26936 19780
rect 31392 19771 31444 19780
rect 28724 19703 28776 19712
rect 28724 19669 28733 19703
rect 28733 19669 28767 19703
rect 28767 19669 28776 19703
rect 28724 19660 28776 19669
rect 29368 19660 29420 19712
rect 31392 19737 31401 19771
rect 31401 19737 31435 19771
rect 31435 19737 31444 19771
rect 31392 19728 31444 19737
rect 41972 19728 42024 19780
rect 31576 19660 31628 19712
rect 34888 19703 34940 19712
rect 34888 19669 34897 19703
rect 34897 19669 34931 19703
rect 34931 19669 34940 19703
rect 34888 19660 34940 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 1768 19456 1820 19508
rect 3792 19456 3844 19508
rect 4528 19456 4580 19508
rect 4896 19456 4948 19508
rect 6092 19456 6144 19508
rect 6276 19456 6328 19508
rect 6644 19456 6696 19508
rect 8944 19456 8996 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 9956 19456 10008 19508
rect 3700 19388 3752 19440
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3608 19320 3660 19372
rect 5816 19388 5868 19440
rect 7472 19388 7524 19440
rect 7564 19388 7616 19440
rect 9128 19388 9180 19440
rect 11060 19388 11112 19440
rect 5632 19320 5684 19372
rect 6276 19320 6328 19372
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 6828 19320 6880 19372
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 10140 19363 10192 19372
rect 10140 19329 10149 19363
rect 10149 19329 10183 19363
rect 10183 19329 10192 19363
rect 10140 19320 10192 19329
rect 11428 19388 11480 19440
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 14004 19456 14056 19508
rect 18328 19499 18380 19508
rect 18328 19465 18337 19499
rect 18337 19465 18371 19499
rect 18371 19465 18380 19499
rect 18328 19456 18380 19465
rect 18512 19456 18564 19508
rect 19248 19456 19300 19508
rect 20628 19456 20680 19508
rect 20812 19456 20864 19508
rect 13728 19388 13780 19440
rect 15016 19388 15068 19440
rect 13820 19320 13872 19372
rect 4528 19295 4580 19304
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 5080 19252 5132 19304
rect 5816 19252 5868 19304
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 10508 19252 10560 19304
rect 12072 19252 12124 19304
rect 12624 19252 12676 19304
rect 14280 19320 14332 19372
rect 14740 19320 14792 19372
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 16580 19320 16632 19372
rect 17316 19320 17368 19372
rect 3332 19227 3384 19236
rect 3332 19193 3341 19227
rect 3341 19193 3375 19227
rect 3375 19193 3384 19227
rect 3332 19184 3384 19193
rect 3792 19116 3844 19168
rect 14004 19252 14056 19304
rect 14096 19252 14148 19304
rect 6276 19116 6328 19168
rect 6920 19116 6972 19168
rect 7564 19116 7616 19168
rect 9128 19116 9180 19168
rect 10784 19116 10836 19168
rect 11152 19116 11204 19168
rect 11428 19116 11480 19168
rect 14188 19184 14240 19236
rect 13084 19116 13136 19168
rect 13544 19116 13596 19168
rect 13728 19116 13780 19168
rect 15016 19116 15068 19168
rect 15200 19116 15252 19168
rect 17224 19252 17276 19304
rect 19340 19388 19392 19440
rect 20260 19388 20312 19440
rect 20536 19388 20588 19440
rect 22468 19499 22520 19508
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 22836 19499 22888 19508
rect 22836 19465 22845 19499
rect 22845 19465 22879 19499
rect 22879 19465 22888 19499
rect 22836 19456 22888 19465
rect 23848 19456 23900 19508
rect 26240 19456 26292 19508
rect 26332 19456 26384 19508
rect 23756 19388 23808 19440
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18604 19320 18656 19372
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 16212 19184 16264 19236
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 20076 19252 20128 19304
rect 20628 19252 20680 19304
rect 20720 19252 20772 19304
rect 21916 19295 21968 19304
rect 21916 19261 21925 19295
rect 21925 19261 21959 19295
rect 21959 19261 21968 19295
rect 21916 19252 21968 19261
rect 25780 19431 25832 19440
rect 25780 19397 25789 19431
rect 25789 19397 25823 19431
rect 25823 19397 25832 19431
rect 25780 19388 25832 19397
rect 25044 19320 25096 19372
rect 16488 19159 16540 19168
rect 16488 19125 16497 19159
rect 16497 19125 16531 19159
rect 16531 19125 16540 19159
rect 16488 19116 16540 19125
rect 16856 19116 16908 19168
rect 18512 19116 18564 19168
rect 22192 19159 22244 19168
rect 22192 19125 22201 19159
rect 22201 19125 22235 19159
rect 22235 19125 22244 19159
rect 22192 19116 22244 19125
rect 23940 19184 23992 19236
rect 28908 19388 28960 19440
rect 29368 19388 29420 19440
rect 26516 19320 26568 19372
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27804 19320 27856 19372
rect 28356 19363 28408 19372
rect 28356 19329 28365 19363
rect 28365 19329 28399 19363
rect 28399 19329 28408 19363
rect 28356 19320 28408 19329
rect 31208 19456 31260 19508
rect 31300 19456 31352 19508
rect 37556 19456 37608 19508
rect 31392 19388 31444 19440
rect 31852 19388 31904 19440
rect 32404 19431 32456 19440
rect 32404 19397 32413 19431
rect 32413 19397 32447 19431
rect 32447 19397 32456 19431
rect 32404 19388 32456 19397
rect 33140 19431 33192 19440
rect 33140 19397 33149 19431
rect 33149 19397 33183 19431
rect 33183 19397 33192 19431
rect 33140 19388 33192 19397
rect 30656 19320 30708 19372
rect 29184 19252 29236 19304
rect 29368 19252 29420 19304
rect 29828 19252 29880 19304
rect 31760 19320 31812 19372
rect 32312 19252 32364 19304
rect 32404 19252 32456 19304
rect 39764 19252 39816 19304
rect 26148 19116 26200 19168
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 45836 19184 45888 19236
rect 32496 19159 32548 19168
rect 32496 19125 32505 19159
rect 32505 19125 32539 19159
rect 32539 19125 32548 19159
rect 32496 19116 32548 19125
rect 33324 19116 33376 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 3424 18912 3476 18964
rect 9128 18912 9180 18964
rect 10416 18912 10468 18964
rect 12440 18912 12492 18964
rect 13728 18912 13780 18964
rect 14464 18912 14516 18964
rect 3608 18887 3660 18896
rect 3608 18853 3617 18887
rect 3617 18853 3651 18887
rect 3651 18853 3660 18887
rect 3608 18844 3660 18853
rect 5080 18844 5132 18896
rect 10600 18887 10652 18896
rect 10600 18853 10609 18887
rect 10609 18853 10643 18887
rect 10643 18853 10652 18887
rect 10600 18844 10652 18853
rect 10968 18844 11020 18896
rect 1400 18776 1452 18828
rect 4160 18776 4212 18828
rect 5356 18776 5408 18828
rect 6828 18776 6880 18828
rect 7380 18776 7432 18828
rect 7840 18776 7892 18828
rect 8576 18776 8628 18828
rect 10140 18776 10192 18828
rect 10324 18776 10376 18828
rect 10692 18776 10744 18828
rect 10876 18776 10928 18828
rect 1860 18708 1912 18760
rect 5264 18640 5316 18692
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 6920 18708 6972 18760
rect 8300 18708 8352 18760
rect 10416 18708 10468 18760
rect 5908 18640 5960 18692
rect 8392 18640 8444 18692
rect 9404 18640 9456 18692
rect 9772 18640 9824 18692
rect 11612 18844 11664 18896
rect 12532 18844 12584 18896
rect 12164 18776 12216 18828
rect 11796 18640 11848 18692
rect 11980 18708 12032 18760
rect 12624 18708 12676 18760
rect 15016 18776 15068 18828
rect 16764 18844 16816 18896
rect 17776 18844 17828 18896
rect 19248 18912 19300 18964
rect 19340 18955 19392 18964
rect 19340 18921 19349 18955
rect 19349 18921 19383 18955
rect 19383 18921 19392 18955
rect 19340 18912 19392 18921
rect 18604 18844 18656 18896
rect 20076 18912 20128 18964
rect 22192 18912 22244 18964
rect 23388 18912 23440 18964
rect 28724 18912 28776 18964
rect 28816 18955 28868 18964
rect 28816 18921 28825 18955
rect 28825 18921 28859 18955
rect 28859 18921 28868 18955
rect 28816 18912 28868 18921
rect 29000 18912 29052 18964
rect 16212 18776 16264 18828
rect 16948 18776 17000 18828
rect 17132 18776 17184 18828
rect 18696 18819 18748 18828
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 14280 18640 14332 18692
rect 15476 18683 15528 18692
rect 15476 18649 15485 18683
rect 15485 18649 15519 18683
rect 15519 18649 15528 18683
rect 15476 18640 15528 18649
rect 16488 18640 16540 18692
rect 7288 18615 7340 18624
rect 7288 18581 7297 18615
rect 7297 18581 7331 18615
rect 7331 18581 7340 18615
rect 7288 18572 7340 18581
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 9036 18572 9088 18624
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 9496 18572 9548 18624
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 11244 18572 11296 18624
rect 11980 18572 12032 18624
rect 12072 18572 12124 18624
rect 12256 18615 12308 18624
rect 12256 18581 12265 18615
rect 12265 18581 12299 18615
rect 12299 18581 12308 18615
rect 12256 18572 12308 18581
rect 17224 18640 17276 18692
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 20168 18776 20220 18828
rect 21456 18819 21508 18828
rect 21456 18785 21465 18819
rect 21465 18785 21499 18819
rect 21499 18785 21508 18819
rect 21456 18776 21508 18785
rect 21824 18776 21876 18828
rect 23940 18776 23992 18828
rect 24032 18776 24084 18828
rect 25780 18776 25832 18828
rect 26148 18776 26200 18828
rect 28448 18844 28500 18896
rect 28632 18887 28684 18896
rect 28632 18853 28641 18887
rect 28641 18853 28675 18887
rect 28675 18853 28684 18887
rect 28632 18844 28684 18853
rect 27252 18776 27304 18828
rect 29828 18776 29880 18828
rect 30012 18776 30064 18828
rect 32404 18844 32456 18896
rect 32588 18844 32640 18896
rect 19708 18708 19760 18760
rect 22468 18708 22520 18760
rect 23296 18708 23348 18760
rect 26792 18708 26844 18760
rect 28632 18708 28684 18760
rect 30196 18751 30248 18760
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 32128 18776 32180 18828
rect 30196 18708 30248 18717
rect 31208 18708 31260 18760
rect 19984 18640 20036 18692
rect 16948 18615 17000 18624
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17408 18572 17460 18624
rect 18236 18572 18288 18624
rect 18512 18572 18564 18624
rect 18604 18615 18656 18624
rect 18604 18581 18613 18615
rect 18613 18581 18647 18615
rect 18647 18581 18656 18615
rect 18604 18572 18656 18581
rect 18696 18572 18748 18624
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 23204 18640 23256 18692
rect 25964 18640 26016 18692
rect 29920 18640 29972 18692
rect 30104 18683 30156 18692
rect 30104 18649 30113 18683
rect 30113 18649 30147 18683
rect 30147 18649 30156 18683
rect 30104 18640 30156 18649
rect 42524 18640 42576 18692
rect 23848 18572 23900 18624
rect 24860 18572 24912 18624
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 25136 18572 25188 18624
rect 27712 18572 27764 18624
rect 29460 18572 29512 18624
rect 29736 18615 29788 18624
rect 29736 18581 29745 18615
rect 29745 18581 29779 18615
rect 29779 18581 29788 18615
rect 29736 18572 29788 18581
rect 30288 18572 30340 18624
rect 32128 18615 32180 18624
rect 32128 18581 32137 18615
rect 32137 18581 32171 18615
rect 32171 18581 32180 18615
rect 32128 18572 32180 18581
rect 43720 18572 43772 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 2228 18368 2280 18420
rect 3792 18300 3844 18352
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 5264 18368 5316 18420
rect 5540 18368 5592 18420
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 14188 18368 14240 18420
rect 15016 18368 15068 18420
rect 17776 18368 17828 18420
rect 6920 18300 6972 18352
rect 8116 18300 8168 18352
rect 9680 18300 9732 18352
rect 9128 18232 9180 18284
rect 9404 18232 9456 18284
rect 11796 18300 11848 18352
rect 14004 18300 14056 18352
rect 19248 18368 19300 18420
rect 12532 18232 12584 18284
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 6000 18164 6052 18216
rect 4896 18096 4948 18148
rect 7288 18164 7340 18216
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 5632 18028 5684 18080
rect 6000 18028 6052 18080
rect 6920 18028 6972 18080
rect 10600 18207 10652 18216
rect 10600 18173 10609 18207
rect 10609 18173 10643 18207
rect 10643 18173 10652 18207
rect 10600 18164 10652 18173
rect 7932 18096 7984 18148
rect 9036 18096 9088 18148
rect 9588 18096 9640 18148
rect 11612 18164 11664 18216
rect 12992 18164 13044 18216
rect 10876 18096 10928 18148
rect 12808 18096 12860 18148
rect 14556 18164 14608 18216
rect 14740 18164 14792 18216
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 17040 18232 17092 18284
rect 20076 18300 20128 18352
rect 13452 18096 13504 18148
rect 11428 18028 11480 18080
rect 12440 18028 12492 18080
rect 13820 18028 13872 18080
rect 14740 18028 14792 18080
rect 16120 18028 16172 18080
rect 16304 18028 16356 18080
rect 16856 18139 16908 18148
rect 16856 18105 16865 18139
rect 16865 18105 16899 18139
rect 16899 18105 16908 18139
rect 16856 18096 16908 18105
rect 18236 18164 18288 18216
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 19984 18232 20036 18284
rect 18972 18164 19024 18216
rect 19616 18096 19668 18148
rect 19800 18164 19852 18216
rect 22652 18368 22704 18420
rect 23204 18368 23256 18420
rect 23388 18368 23440 18420
rect 25044 18368 25096 18420
rect 20352 18207 20404 18216
rect 20352 18173 20361 18207
rect 20361 18173 20395 18207
rect 20395 18173 20404 18207
rect 20352 18164 20404 18173
rect 23664 18300 23716 18352
rect 27712 18368 27764 18420
rect 25964 18300 26016 18352
rect 29368 18368 29420 18420
rect 29828 18411 29880 18420
rect 29828 18377 29837 18411
rect 29837 18377 29871 18411
rect 29871 18377 29880 18411
rect 29828 18368 29880 18377
rect 37188 18368 37240 18420
rect 28356 18300 28408 18352
rect 29644 18300 29696 18352
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 19340 18071 19392 18080
rect 19340 18037 19349 18071
rect 19349 18037 19383 18071
rect 19383 18037 19392 18071
rect 19340 18028 19392 18037
rect 19432 18028 19484 18080
rect 20352 18028 20404 18080
rect 20444 18028 20496 18080
rect 20904 18028 20956 18080
rect 21364 18028 21416 18080
rect 24400 18232 24452 18284
rect 26792 18232 26844 18284
rect 28080 18275 28132 18284
rect 28080 18241 28089 18275
rect 28089 18241 28123 18275
rect 28123 18241 28132 18275
rect 28080 18232 28132 18241
rect 29460 18232 29512 18284
rect 31116 18232 31168 18284
rect 23756 18164 23808 18216
rect 30288 18164 30340 18216
rect 30840 18207 30892 18216
rect 30840 18173 30849 18207
rect 30849 18173 30883 18207
rect 30883 18173 30892 18207
rect 30840 18164 30892 18173
rect 24768 18096 24820 18148
rect 31760 18139 31812 18148
rect 31760 18105 31769 18139
rect 31769 18105 31803 18139
rect 31803 18105 31812 18139
rect 31760 18096 31812 18105
rect 25320 18028 25372 18080
rect 26516 18028 26568 18080
rect 26792 18028 26844 18080
rect 27436 18028 27488 18080
rect 29460 18028 29512 18080
rect 30288 18071 30340 18080
rect 30288 18037 30297 18071
rect 30297 18037 30331 18071
rect 30331 18037 30340 18071
rect 30288 18028 30340 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 6184 17824 6236 17876
rect 10324 17824 10376 17876
rect 10508 17824 10560 17876
rect 1216 17688 1268 17740
rect 6736 17756 6788 17808
rect 3884 17688 3936 17740
rect 4620 17688 4672 17740
rect 6552 17688 6604 17740
rect 8116 17688 8168 17740
rect 13820 17824 13872 17876
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 14832 17867 14884 17876
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 15844 17824 15896 17876
rect 14004 17756 14056 17808
rect 15200 17756 15252 17808
rect 19248 17824 19300 17876
rect 20444 17756 20496 17808
rect 20904 17756 20956 17808
rect 11336 17688 11388 17740
rect 11612 17688 11664 17740
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 14556 17688 14608 17740
rect 16212 17688 16264 17740
rect 20628 17688 20680 17740
rect 20812 17688 20864 17740
rect 21732 17867 21784 17876
rect 21732 17833 21741 17867
rect 21741 17833 21775 17867
rect 21775 17833 21784 17867
rect 21732 17824 21784 17833
rect 21916 17867 21968 17876
rect 21916 17833 21925 17867
rect 21925 17833 21959 17867
rect 21959 17833 21968 17867
rect 21916 17824 21968 17833
rect 24032 17824 24084 17876
rect 24768 17824 24820 17876
rect 26516 17824 26568 17876
rect 27620 17824 27672 17876
rect 28908 17867 28960 17876
rect 28908 17833 28917 17867
rect 28917 17833 28951 17867
rect 28951 17833 28960 17867
rect 28908 17824 28960 17833
rect 30840 17824 30892 17876
rect 31116 17824 31168 17876
rect 30380 17756 30432 17808
rect 32496 17756 32548 17808
rect 23756 17688 23808 17740
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 7012 17620 7064 17672
rect 1400 17552 1452 17604
rect 4804 17552 4856 17604
rect 6644 17552 6696 17604
rect 6828 17552 6880 17604
rect 3884 17484 3936 17536
rect 6552 17484 6604 17536
rect 7104 17484 7156 17536
rect 8208 17484 8260 17536
rect 9128 17595 9180 17604
rect 9128 17561 9137 17595
rect 9137 17561 9171 17595
rect 9171 17561 9180 17595
rect 9128 17552 9180 17561
rect 9864 17595 9916 17604
rect 9864 17561 9873 17595
rect 9873 17561 9907 17595
rect 9907 17561 9916 17595
rect 9864 17552 9916 17561
rect 9680 17484 9732 17536
rect 10600 17484 10652 17536
rect 10784 17484 10836 17536
rect 13636 17620 13688 17672
rect 15844 17620 15896 17672
rect 19432 17620 19484 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 20076 17620 20128 17672
rect 11336 17552 11388 17604
rect 12440 17552 12492 17604
rect 13820 17552 13872 17604
rect 13912 17552 13964 17604
rect 16488 17552 16540 17604
rect 20168 17552 20220 17604
rect 20260 17595 20312 17604
rect 20260 17561 20269 17595
rect 20269 17561 20303 17595
rect 20303 17561 20312 17595
rect 20260 17552 20312 17561
rect 14096 17484 14148 17536
rect 14280 17484 14332 17536
rect 14464 17484 14516 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 17224 17484 17276 17536
rect 21088 17620 21140 17672
rect 21640 17552 21692 17604
rect 23848 17552 23900 17604
rect 24308 17552 24360 17604
rect 21364 17484 21416 17536
rect 21824 17484 21876 17536
rect 21916 17484 21968 17536
rect 22468 17484 22520 17536
rect 23296 17484 23348 17536
rect 24124 17484 24176 17536
rect 24952 17731 25004 17740
rect 24952 17697 24961 17731
rect 24961 17697 24995 17731
rect 24995 17697 25004 17731
rect 24952 17688 25004 17697
rect 27804 17688 27856 17740
rect 28080 17688 28132 17740
rect 28724 17688 28776 17740
rect 29460 17620 29512 17672
rect 30012 17688 30064 17740
rect 31300 17688 31352 17740
rect 31024 17620 31076 17672
rect 24860 17552 24912 17604
rect 26792 17552 26844 17604
rect 27712 17552 27764 17604
rect 45468 17552 45520 17604
rect 29368 17484 29420 17536
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 47032 17484 47084 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 5540 17280 5592 17332
rect 9220 17280 9272 17332
rect 9404 17280 9456 17332
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 10324 17280 10376 17332
rect 4252 17212 4304 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 13360 17212 13412 17264
rect 20260 17280 20312 17332
rect 21272 17280 21324 17332
rect 30288 17280 30340 17332
rect 14188 17212 14240 17264
rect 15568 17212 15620 17264
rect 15844 17212 15896 17264
rect 21824 17255 21876 17264
rect 21824 17221 21833 17255
rect 21833 17221 21867 17255
rect 21867 17221 21876 17255
rect 21824 17212 21876 17221
rect 23480 17212 23532 17264
rect 23940 17255 23992 17264
rect 23940 17221 23949 17255
rect 23949 17221 23983 17255
rect 23983 17221 23992 17255
rect 23940 17212 23992 17221
rect 24032 17255 24084 17264
rect 24032 17221 24041 17255
rect 24041 17221 24075 17255
rect 24075 17221 24084 17255
rect 24032 17212 24084 17221
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 1308 17076 1360 17128
rect 2872 17076 2924 17128
rect 6644 17144 6696 17196
rect 4896 17008 4948 17060
rect 6368 17008 6420 17060
rect 5540 16940 5592 16992
rect 6184 16940 6236 16992
rect 8392 17187 8444 17196
rect 8392 17153 8401 17187
rect 8401 17153 8435 17187
rect 8435 17153 8444 17187
rect 8392 17144 8444 17153
rect 7288 17008 7340 17060
rect 9956 17144 10008 17196
rect 8852 17076 8904 17128
rect 9036 17076 9088 17128
rect 10232 17076 10284 17128
rect 10324 17076 10376 17128
rect 10692 17008 10744 17060
rect 7932 16940 7984 16992
rect 8208 16940 8260 16992
rect 8300 16940 8352 16992
rect 9772 16940 9824 16992
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 10876 16940 10928 16992
rect 11428 17144 11480 17196
rect 12072 17144 12124 17196
rect 12624 17076 12676 17128
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 14096 17144 14148 17196
rect 14280 17144 14332 17196
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 16672 17144 16724 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 24952 17212 25004 17264
rect 26792 17212 26844 17264
rect 29460 17212 29512 17264
rect 31300 17212 31352 17264
rect 12440 17051 12492 17060
rect 12440 17017 12449 17051
rect 12449 17017 12483 17051
rect 12483 17017 12492 17051
rect 12440 17008 12492 17017
rect 12532 17008 12584 17060
rect 15936 17076 15988 17128
rect 17776 17076 17828 17128
rect 13728 17008 13780 17060
rect 16764 17008 16816 17060
rect 17132 17008 17184 17060
rect 19616 17076 19668 17128
rect 27804 17144 27856 17196
rect 19800 17008 19852 17060
rect 11796 16940 11848 16992
rect 13452 16940 13504 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 14004 16940 14056 16992
rect 15384 16940 15436 16992
rect 16580 16940 16632 16992
rect 17040 16940 17092 16992
rect 20076 16940 20128 16992
rect 20628 16940 20680 16992
rect 20904 16940 20956 16992
rect 21180 17008 21232 17060
rect 21732 16940 21784 16992
rect 21916 16940 21968 16992
rect 23480 16940 23532 16992
rect 23572 16983 23624 16992
rect 23572 16949 23581 16983
rect 23581 16949 23615 16983
rect 23615 16949 23624 16983
rect 23572 16940 23624 16949
rect 23940 17076 23992 17128
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 30012 17076 30064 17128
rect 26148 17008 26200 17060
rect 32864 17008 32916 17060
rect 34520 17008 34572 17060
rect 27528 16940 27580 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 5080 16736 5132 16788
rect 6092 16736 6144 16788
rect 2228 16600 2280 16652
rect 9680 16736 9732 16788
rect 12072 16736 12124 16788
rect 12256 16736 12308 16788
rect 3332 16600 3384 16652
rect 7104 16643 7156 16652
rect 7104 16609 7113 16643
rect 7113 16609 7147 16643
rect 7147 16609 7156 16643
rect 7104 16600 7156 16609
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 1308 16464 1360 16516
rect 4712 16532 4764 16584
rect 7840 16532 7892 16584
rect 8116 16600 8168 16652
rect 8668 16668 8720 16720
rect 9404 16668 9456 16720
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 8760 16532 8812 16584
rect 10600 16532 10652 16584
rect 11796 16532 11848 16584
rect 12072 16532 12124 16584
rect 14188 16736 14240 16788
rect 14464 16779 14516 16788
rect 14464 16745 14473 16779
rect 14473 16745 14507 16779
rect 14507 16745 14516 16779
rect 14464 16736 14516 16745
rect 14648 16736 14700 16788
rect 18972 16736 19024 16788
rect 20076 16736 20128 16788
rect 23020 16736 23072 16788
rect 23296 16779 23348 16788
rect 23296 16745 23305 16779
rect 23305 16745 23339 16779
rect 23339 16745 23348 16779
rect 23296 16736 23348 16745
rect 24124 16736 24176 16788
rect 16948 16668 17000 16720
rect 18512 16668 18564 16720
rect 18880 16668 18932 16720
rect 20720 16668 20772 16720
rect 12624 16600 12676 16652
rect 13268 16600 13320 16652
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 14372 16600 14424 16652
rect 15016 16532 15068 16584
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16304 16600 16356 16652
rect 6276 16464 6328 16516
rect 7104 16464 7156 16516
rect 8576 16464 8628 16516
rect 9864 16464 9916 16516
rect 10140 16464 10192 16516
rect 11428 16464 11480 16516
rect 12440 16464 12492 16516
rect 13544 16464 13596 16516
rect 14648 16464 14700 16516
rect 15752 16464 15804 16516
rect 16212 16532 16264 16584
rect 16764 16532 16816 16584
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18604 16600 18656 16652
rect 19156 16600 19208 16652
rect 21088 16600 21140 16652
rect 21824 16600 21876 16652
rect 21916 16600 21968 16652
rect 19248 16532 19300 16584
rect 19800 16464 19852 16516
rect 20444 16464 20496 16516
rect 21272 16464 21324 16516
rect 5448 16396 5500 16448
rect 6460 16396 6512 16448
rect 7564 16396 7616 16448
rect 7656 16396 7708 16448
rect 9220 16396 9272 16448
rect 11060 16396 11112 16448
rect 12624 16396 12676 16448
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 17408 16396 17460 16448
rect 18420 16439 18472 16448
rect 18420 16405 18429 16439
rect 18429 16405 18463 16439
rect 18463 16405 18472 16439
rect 18420 16396 18472 16405
rect 19064 16396 19116 16448
rect 22284 16532 22336 16584
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 24952 16600 25004 16652
rect 25688 16600 25740 16652
rect 26056 16600 26108 16652
rect 29736 16668 29788 16720
rect 27804 16643 27856 16652
rect 27804 16609 27813 16643
rect 27813 16609 27847 16643
rect 27847 16609 27856 16643
rect 27804 16600 27856 16609
rect 28724 16600 28776 16652
rect 31484 16668 31536 16720
rect 30012 16643 30064 16652
rect 30012 16609 30021 16643
rect 30021 16609 30055 16643
rect 30055 16609 30064 16643
rect 30012 16600 30064 16609
rect 23756 16532 23808 16584
rect 23020 16507 23072 16516
rect 23020 16473 23029 16507
rect 23029 16473 23063 16507
rect 23063 16473 23072 16507
rect 26424 16532 26476 16584
rect 27252 16532 27304 16584
rect 29552 16532 29604 16584
rect 23020 16464 23072 16473
rect 25320 16464 25372 16516
rect 22192 16396 22244 16448
rect 22652 16396 22704 16448
rect 23204 16396 23256 16448
rect 23664 16396 23716 16448
rect 24768 16439 24820 16448
rect 24768 16405 24777 16439
rect 24777 16405 24811 16439
rect 24811 16405 24820 16439
rect 24768 16396 24820 16405
rect 27252 16439 27304 16448
rect 27252 16405 27261 16439
rect 27261 16405 27295 16439
rect 27295 16405 27304 16439
rect 27252 16396 27304 16405
rect 29368 16464 29420 16516
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 480 16192 532 16244
rect 1124 16192 1176 16244
rect 3792 16192 3844 16244
rect 4436 16167 4488 16176
rect 4436 16133 4445 16167
rect 4445 16133 4479 16167
rect 4479 16133 4488 16167
rect 4436 16124 4488 16133
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 6552 16192 6604 16244
rect 8668 16192 8720 16244
rect 8852 16192 8904 16244
rect 8944 16235 8996 16244
rect 8944 16201 8953 16235
rect 8953 16201 8987 16235
rect 8987 16201 8996 16235
rect 8944 16192 8996 16201
rect 9404 16192 9456 16244
rect 16488 16192 16540 16244
rect 17040 16192 17092 16244
rect 3332 16056 3384 16108
rect 1308 15988 1360 16040
rect 4804 15988 4856 16040
rect 6368 15988 6420 16040
rect 7012 16099 7064 16108
rect 7012 16065 7021 16099
rect 7021 16065 7055 16099
rect 7055 16065 7064 16099
rect 7012 16056 7064 16065
rect 8392 16124 8444 16176
rect 8576 16056 8628 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 7656 15988 7708 16040
rect 7748 15988 7800 16040
rect 8668 15988 8720 16040
rect 9404 16056 9456 16108
rect 10140 16056 10192 16108
rect 10508 16167 10560 16176
rect 10508 16133 10517 16167
rect 10517 16133 10551 16167
rect 10551 16133 10560 16167
rect 10508 16124 10560 16133
rect 12256 16124 12308 16176
rect 13820 16124 13872 16176
rect 14096 16124 14148 16176
rect 14372 16124 14424 16176
rect 19064 16192 19116 16244
rect 10876 16056 10928 16108
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 13268 16056 13320 16108
rect 14648 16056 14700 16108
rect 15292 16056 15344 16108
rect 7932 15920 7984 15972
rect 8484 15963 8536 15972
rect 8484 15929 8493 15963
rect 8493 15929 8527 15963
rect 8527 15929 8536 15963
rect 8484 15920 8536 15929
rect 6552 15852 6604 15904
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 8576 15852 8628 15904
rect 10600 16031 10652 16040
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 10692 16031 10744 16040
rect 10692 15997 10701 16031
rect 10701 15997 10735 16031
rect 10735 15997 10744 16031
rect 10692 15988 10744 15997
rect 12992 15988 13044 16040
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 16028 16056 16080 16108
rect 19432 16124 19484 16176
rect 20536 16124 20588 16176
rect 23296 16192 23348 16244
rect 27252 16192 27304 16244
rect 26424 16124 26476 16176
rect 27804 16124 27856 16176
rect 43536 16124 43588 16176
rect 19064 16056 19116 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 21548 16056 21600 16108
rect 23572 16056 23624 16108
rect 26516 16056 26568 16108
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27528 16056 27580 16108
rect 28908 16056 28960 16108
rect 18604 15988 18656 16040
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 22468 15988 22520 16040
rect 13636 15920 13688 15972
rect 15660 15920 15712 15972
rect 18512 15920 18564 15972
rect 18788 15920 18840 15972
rect 18972 15920 19024 15972
rect 20168 15920 20220 15972
rect 9496 15852 9548 15904
rect 9864 15852 9916 15904
rect 10600 15852 10652 15904
rect 11060 15852 11112 15904
rect 11612 15852 11664 15904
rect 11796 15852 11848 15904
rect 11980 15852 12032 15904
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 16028 15852 16080 15904
rect 16488 15852 16540 15904
rect 17316 15852 17368 15904
rect 19616 15895 19668 15904
rect 19616 15861 19625 15895
rect 19625 15861 19659 15895
rect 19659 15861 19668 15895
rect 19616 15852 19668 15861
rect 20720 15852 20772 15904
rect 21732 15852 21784 15904
rect 23204 15988 23256 16040
rect 22744 15920 22796 15972
rect 23572 15852 23624 15904
rect 24860 16031 24912 16040
rect 24860 15997 24869 16031
rect 24869 15997 24903 16031
rect 24903 15997 24912 16031
rect 24860 15988 24912 15997
rect 26148 15920 26200 15972
rect 27620 15852 27672 15904
rect 27712 15852 27764 15904
rect 29552 15895 29604 15904
rect 29552 15861 29561 15895
rect 29561 15861 29595 15895
rect 29595 15861 29604 15895
rect 29552 15852 29604 15861
rect 30380 15920 30432 15972
rect 46940 15920 46992 15972
rect 45284 15852 45336 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 5632 15648 5684 15700
rect 6736 15580 6788 15632
rect 7564 15648 7616 15700
rect 7932 15648 7984 15700
rect 9404 15648 9456 15700
rect 9634 15648 9686 15700
rect 10508 15648 10560 15700
rect 10600 15648 10652 15700
rect 1308 15512 1360 15564
rect 4896 15512 4948 15564
rect 6368 15512 6420 15564
rect 6552 15512 6604 15564
rect 8760 15580 8812 15632
rect 8484 15555 8536 15564
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 8484 15512 8536 15521
rect 8668 15512 8720 15564
rect 9772 15580 9824 15632
rect 11428 15580 11480 15632
rect 13452 15648 13504 15700
rect 15476 15648 15528 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 17776 15648 17828 15700
rect 18972 15648 19024 15700
rect 9634 15512 9686 15564
rect 10324 15555 10376 15564
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 10600 15512 10652 15564
rect 3516 15444 3568 15496
rect 4252 15444 4304 15496
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 7840 15444 7892 15496
rect 7932 15444 7984 15496
rect 9864 15444 9916 15496
rect 10416 15444 10468 15496
rect 11612 15444 11664 15496
rect 2688 15308 2740 15360
rect 3792 15308 3844 15360
rect 6460 15376 6512 15428
rect 8668 15376 8720 15428
rect 9404 15376 9456 15428
rect 9588 15376 9640 15428
rect 11428 15419 11480 15428
rect 11428 15385 11437 15419
rect 11437 15385 11471 15419
rect 11471 15385 11480 15419
rect 11428 15376 11480 15385
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 5448 15308 5500 15360
rect 7472 15308 7524 15360
rect 8760 15308 8812 15360
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 9864 15308 9916 15360
rect 11520 15308 11572 15360
rect 13636 15512 13688 15564
rect 14832 15512 14884 15564
rect 15660 15512 15712 15564
rect 16764 15512 16816 15564
rect 13268 15444 13320 15496
rect 15568 15444 15620 15496
rect 16856 15444 16908 15496
rect 15200 15376 15252 15428
rect 16764 15376 16816 15428
rect 12164 15351 12216 15360
rect 12164 15317 12173 15351
rect 12173 15317 12207 15351
rect 12207 15317 12216 15351
rect 12164 15308 12216 15317
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 16212 15308 16264 15360
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 20536 15580 20588 15632
rect 22468 15580 22520 15632
rect 19432 15512 19484 15564
rect 20168 15555 20220 15564
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 20996 15512 21048 15564
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 22100 15512 22152 15564
rect 23848 15555 23900 15564
rect 23848 15521 23857 15555
rect 23857 15521 23891 15555
rect 23891 15521 23900 15555
rect 23848 15512 23900 15521
rect 26608 15648 26660 15700
rect 24952 15580 25004 15632
rect 25688 15512 25740 15564
rect 26884 15555 26936 15564
rect 26884 15521 26893 15555
rect 26893 15521 26927 15555
rect 26927 15521 26936 15555
rect 26884 15512 26936 15521
rect 28540 15648 28592 15700
rect 28724 15648 28776 15700
rect 27160 15444 27212 15496
rect 27620 15487 27672 15496
rect 27620 15453 27629 15487
rect 27629 15453 27663 15487
rect 27663 15453 27672 15487
rect 27620 15444 27672 15453
rect 17408 15419 17460 15428
rect 17408 15385 17417 15419
rect 17417 15385 17451 15419
rect 17451 15385 17460 15419
rect 17408 15376 17460 15385
rect 18972 15376 19024 15428
rect 18880 15308 18932 15360
rect 19248 15308 19300 15360
rect 20076 15351 20128 15360
rect 20076 15317 20085 15351
rect 20085 15317 20119 15351
rect 20119 15317 20128 15351
rect 20076 15308 20128 15317
rect 20628 15376 20680 15428
rect 21088 15376 21140 15428
rect 21364 15419 21416 15428
rect 21364 15385 21373 15419
rect 21373 15385 21407 15419
rect 21407 15385 21416 15419
rect 21364 15376 21416 15385
rect 23572 15376 23624 15428
rect 23664 15419 23716 15428
rect 23664 15385 23673 15419
rect 23673 15385 23707 15419
rect 23707 15385 23716 15419
rect 23664 15376 23716 15385
rect 24308 15376 24360 15428
rect 26148 15376 26200 15428
rect 27804 15376 27856 15428
rect 21732 15308 21784 15360
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 24400 15308 24452 15360
rect 25228 15351 25280 15360
rect 25228 15317 25237 15351
rect 25237 15317 25271 15351
rect 25271 15317 25280 15351
rect 25228 15308 25280 15317
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 25780 15308 25832 15360
rect 26976 15308 27028 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 204 15104 256 15156
rect 1124 15104 1176 15156
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 4988 15147 5040 15156
rect 4988 15113 4997 15147
rect 4997 15113 5031 15147
rect 5031 15113 5040 15147
rect 4988 15104 5040 15113
rect 6552 15104 6604 15156
rect 7840 15104 7892 15156
rect 8208 15104 8260 15156
rect 8484 15104 8536 15156
rect 3424 14968 3476 15020
rect 8760 15036 8812 15088
rect 9496 15036 9548 15088
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 6184 14968 6236 15020
rect 6368 14968 6420 15020
rect 1124 14900 1176 14952
rect 4160 14900 4212 14952
rect 5632 14900 5684 14952
rect 6920 14968 6972 15020
rect 9956 15079 10008 15088
rect 9956 15045 9965 15079
rect 9965 15045 9999 15079
rect 9999 15045 10008 15079
rect 9956 15036 10008 15045
rect 10140 15036 10192 15088
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 18236 15104 18288 15156
rect 19524 15104 19576 15156
rect 20628 15104 20680 15156
rect 20720 15104 20772 15156
rect 21272 15104 21324 15156
rect 21364 15104 21416 15156
rect 27160 15104 27212 15156
rect 27436 15147 27488 15156
rect 27436 15113 27445 15147
rect 27445 15113 27479 15147
rect 27479 15113 27488 15147
rect 27436 15104 27488 15113
rect 27804 15104 27856 15156
rect 10692 14968 10744 15020
rect 7748 14900 7800 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 10600 14900 10652 14952
rect 11612 14968 11664 15020
rect 13268 15036 13320 15088
rect 16396 15036 16448 15088
rect 19340 15036 19392 15088
rect 19616 15036 19668 15088
rect 20536 15036 20588 15088
rect 22100 15036 22152 15088
rect 24860 15036 24912 15088
rect 26884 15036 26936 15088
rect 12808 15011 12860 15020
rect 12808 14977 12817 15011
rect 12817 14977 12851 15011
rect 12851 14977 12860 15011
rect 12808 14968 12860 14977
rect 13544 14968 13596 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 16304 14968 16356 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 19432 14968 19484 15020
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 13728 14900 13780 14952
rect 16212 14900 16264 14952
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 8944 14764 8996 14816
rect 9588 14764 9640 14816
rect 9956 14764 10008 14816
rect 10508 14764 10560 14816
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 16948 14900 17000 14952
rect 17408 14900 17460 14952
rect 20720 14900 20772 14952
rect 20996 14900 21048 14952
rect 22468 14968 22520 15020
rect 23388 14968 23440 15020
rect 26516 14968 26568 15020
rect 27436 14968 27488 15020
rect 27620 14968 27672 15020
rect 16764 14832 16816 14884
rect 18236 14832 18288 14884
rect 18788 14832 18840 14884
rect 19156 14832 19208 14884
rect 13544 14764 13596 14773
rect 16948 14764 17000 14816
rect 19340 14764 19392 14816
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 21364 14832 21416 14884
rect 20996 14764 21048 14816
rect 22560 14764 22612 14816
rect 24308 14807 24360 14816
rect 24308 14773 24317 14807
rect 24317 14773 24351 14807
rect 24351 14773 24360 14807
rect 24308 14764 24360 14773
rect 24400 14764 24452 14816
rect 24860 14764 24912 14816
rect 26976 14900 27028 14952
rect 26148 14832 26200 14884
rect 43444 14900 43496 14952
rect 25872 14764 25924 14816
rect 26240 14764 26292 14816
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 27436 14764 27488 14816
rect 46204 14832 46256 14884
rect 48596 14764 48648 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 4160 14603 4212 14612
rect 4160 14569 4169 14603
rect 4169 14569 4203 14603
rect 4203 14569 4212 14603
rect 4160 14560 4212 14569
rect 8484 14560 8536 14612
rect 1308 14424 1360 14476
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 4804 14467 4856 14476
rect 4804 14433 4813 14467
rect 4813 14433 4847 14467
rect 4847 14433 4856 14467
rect 4804 14424 4856 14433
rect 4896 14424 4948 14476
rect 7656 14492 7708 14544
rect 7564 14424 7616 14476
rect 8208 14424 8260 14476
rect 9220 14492 9272 14544
rect 5172 14356 5224 14408
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 8484 14424 8536 14476
rect 9772 14492 9824 14544
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 14096 14560 14148 14612
rect 11980 14492 12032 14544
rect 13544 14492 13596 14544
rect 17316 14560 17368 14612
rect 18512 14560 18564 14612
rect 18696 14560 18748 14612
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 10140 14424 10192 14476
rect 10232 14424 10284 14476
rect 10600 14356 10652 14408
rect 10876 14356 10928 14408
rect 14188 14424 14240 14476
rect 15384 14424 15436 14476
rect 18420 14424 18472 14476
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 19248 14560 19300 14612
rect 19984 14560 20036 14612
rect 20628 14560 20680 14612
rect 21824 14560 21876 14612
rect 25688 14560 25740 14612
rect 27160 14603 27212 14612
rect 27160 14569 27169 14603
rect 27169 14569 27203 14603
rect 27203 14569 27212 14603
rect 27160 14560 27212 14569
rect 24860 14492 24912 14544
rect 26332 14492 26384 14544
rect 19340 14424 19392 14476
rect 20168 14424 20220 14476
rect 22100 14424 22152 14476
rect 4160 14288 4212 14340
rect 5540 14288 5592 14340
rect 7748 14288 7800 14340
rect 3332 14263 3384 14272
rect 3332 14229 3341 14263
rect 3341 14229 3375 14263
rect 3375 14229 3384 14263
rect 3332 14220 3384 14229
rect 4436 14220 4488 14272
rect 4804 14220 4856 14272
rect 7288 14220 7340 14272
rect 8484 14220 8536 14272
rect 8852 14220 8904 14272
rect 9588 14220 9640 14272
rect 9864 14220 9916 14272
rect 11060 14220 11112 14272
rect 11704 14220 11756 14272
rect 12532 14288 12584 14340
rect 13728 14288 13780 14340
rect 16304 14288 16356 14340
rect 15936 14220 15988 14272
rect 21364 14356 21416 14408
rect 23664 14356 23716 14408
rect 23940 14356 23992 14408
rect 17040 14288 17092 14340
rect 18696 14288 18748 14340
rect 17132 14220 17184 14272
rect 19064 14220 19116 14272
rect 19984 14220 20036 14272
rect 20996 14331 21048 14340
rect 20996 14297 21005 14331
rect 21005 14297 21039 14331
rect 21039 14297 21048 14331
rect 20996 14288 21048 14297
rect 21180 14288 21232 14340
rect 21824 14288 21876 14340
rect 22468 14288 22520 14340
rect 22560 14331 22612 14340
rect 22560 14297 22569 14331
rect 22569 14297 22603 14331
rect 22603 14297 22612 14331
rect 22560 14288 22612 14297
rect 20904 14220 20956 14272
rect 25964 14331 26016 14340
rect 25964 14297 25973 14331
rect 25973 14297 26007 14331
rect 26007 14297 26016 14331
rect 25964 14288 26016 14297
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 24952 14220 25004 14272
rect 26516 14220 26568 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 112 13880 164 13932
rect 756 13880 808 13932
rect 3608 13880 3660 13932
rect 5816 14016 5868 14068
rect 6460 14059 6512 14068
rect 6460 14025 6469 14059
rect 6469 14025 6503 14059
rect 6503 14025 6512 14059
rect 6460 14016 6512 14025
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7840 14016 7892 14068
rect 8300 14016 8352 14068
rect 8576 14059 8628 14068
rect 8576 14025 8585 14059
rect 8585 14025 8619 14059
rect 8619 14025 8628 14059
rect 8576 14016 8628 14025
rect 8944 14016 8996 14068
rect 10232 14016 10284 14068
rect 10324 14016 10376 14068
rect 11612 14016 11664 14068
rect 12900 14016 12952 14068
rect 13268 14016 13320 14068
rect 13360 14059 13412 14068
rect 13360 14025 13369 14059
rect 13369 14025 13403 14059
rect 13403 14025 13412 14059
rect 13360 14016 13412 14025
rect 15292 14016 15344 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 17224 14016 17276 14068
rect 5080 13948 5132 14000
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 5540 13880 5592 13932
rect 1308 13812 1360 13864
rect 4988 13812 5040 13864
rect 5080 13812 5132 13864
rect 5632 13812 5684 13864
rect 6184 13812 6236 13864
rect 6368 13812 6420 13864
rect 6644 13948 6696 14000
rect 8760 13948 8812 14000
rect 9496 13948 9548 14000
rect 7748 13880 7800 13932
rect 13544 13948 13596 14000
rect 13820 13948 13872 14000
rect 16304 13948 16356 14000
rect 17040 13948 17092 14000
rect 17868 13948 17920 14000
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 19248 14059 19300 14068
rect 19248 14025 19257 14059
rect 19257 14025 19291 14059
rect 19291 14025 19300 14059
rect 19248 14016 19300 14025
rect 20444 14016 20496 14068
rect 20628 14016 20680 14068
rect 20996 14016 21048 14068
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 20720 13948 20772 14000
rect 24124 14016 24176 14068
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 26148 14016 26200 14068
rect 26332 14016 26384 14068
rect 27712 14016 27764 14068
rect 24860 13948 24912 14000
rect 25596 13948 25648 14000
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 6828 13812 6880 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 756 13744 808 13796
rect 1216 13744 1268 13796
rect 3792 13676 3844 13728
rect 8484 13744 8536 13796
rect 12164 13880 12216 13932
rect 15660 13880 15712 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 20536 13923 20588 13932
rect 20536 13889 20545 13923
rect 20545 13889 20579 13923
rect 20579 13889 20588 13923
rect 20536 13880 20588 13889
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 9588 13855 9640 13864
rect 9588 13821 9597 13855
rect 9597 13821 9631 13855
rect 9631 13821 9640 13855
rect 9588 13812 9640 13821
rect 10232 13812 10284 13864
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 10968 13744 11020 13796
rect 12348 13744 12400 13796
rect 9588 13676 9640 13728
rect 10324 13676 10376 13728
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13728 13812 13780 13864
rect 15384 13812 15436 13864
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 12716 13744 12768 13796
rect 13820 13787 13872 13796
rect 13820 13753 13829 13787
rect 13829 13753 13863 13787
rect 13863 13753 13872 13787
rect 13820 13744 13872 13753
rect 14372 13744 14424 13796
rect 16488 13744 16540 13796
rect 17500 13812 17552 13864
rect 18512 13744 18564 13796
rect 18972 13744 19024 13796
rect 20904 13812 20956 13864
rect 22192 13880 22244 13932
rect 23480 13880 23532 13932
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 24584 13880 24636 13889
rect 21824 13744 21876 13796
rect 22652 13744 22704 13796
rect 24308 13812 24360 13864
rect 30380 13880 30432 13932
rect 24492 13744 24544 13796
rect 24952 13744 25004 13796
rect 26240 13744 26292 13796
rect 15660 13676 15712 13728
rect 17960 13676 18012 13728
rect 22100 13676 22152 13728
rect 23940 13676 23992 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 6000 13472 6052 13524
rect 3424 13447 3476 13456
rect 3424 13413 3433 13447
rect 3433 13413 3467 13447
rect 3467 13413 3476 13447
rect 3424 13404 3476 13413
rect 3884 13404 3936 13456
rect 5080 13404 5132 13456
rect 5264 13404 5316 13456
rect 7196 13472 7248 13524
rect 7472 13472 7524 13524
rect 15108 13472 15160 13524
rect 17592 13472 17644 13524
rect 20720 13472 20772 13524
rect 22100 13472 22152 13524
rect 22468 13472 22520 13524
rect 23388 13472 23440 13524
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 4620 13336 4672 13388
rect 6000 13336 6052 13388
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 7564 13336 7616 13388
rect 7748 13336 7800 13388
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 11060 13404 11112 13456
rect 11704 13404 11756 13456
rect 13636 13404 13688 13456
rect 15660 13404 15712 13456
rect 16856 13404 16908 13456
rect 18604 13404 18656 13456
rect 24308 13404 24360 13456
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 3884 13268 3936 13320
rect 4344 13268 4396 13320
rect 5448 13268 5500 13320
rect 5816 13268 5868 13320
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8484 13268 8536 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 12256 13336 12308 13388
rect 14648 13336 14700 13388
rect 15108 13336 15160 13388
rect 16672 13336 16724 13388
rect 17132 13379 17184 13388
rect 17132 13345 17141 13379
rect 17141 13345 17175 13379
rect 17175 13345 17184 13379
rect 17132 13336 17184 13345
rect 19708 13336 19760 13388
rect 20904 13336 20956 13388
rect 22192 13336 22244 13388
rect 11336 13268 11388 13320
rect 16028 13268 16080 13320
rect 16948 13268 17000 13320
rect 18420 13268 18472 13320
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 21916 13268 21968 13320
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 23940 13336 23992 13388
rect 24400 13268 24452 13320
rect 25044 13268 25096 13320
rect 25688 13268 25740 13320
rect 6276 13200 6328 13252
rect 7196 13200 7248 13252
rect 4436 13132 4488 13184
rect 5724 13132 5776 13184
rect 5816 13132 5868 13184
rect 9220 13132 9272 13184
rect 9404 13132 9456 13184
rect 10140 13132 10192 13184
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 11704 13200 11756 13252
rect 13728 13200 13780 13252
rect 14004 13132 14056 13184
rect 16672 13200 16724 13252
rect 18052 13200 18104 13252
rect 21088 13200 21140 13252
rect 15936 13132 15988 13184
rect 17316 13132 17368 13184
rect 17776 13132 17828 13184
rect 18328 13132 18380 13184
rect 32220 13200 32272 13252
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 23664 13132 23716 13184
rect 24492 13132 24544 13184
rect 25780 13132 25832 13184
rect 26424 13175 26476 13184
rect 26424 13141 26433 13175
rect 26433 13141 26467 13175
rect 26467 13141 26476 13175
rect 26424 13132 26476 13141
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3332 12928 3384 12980
rect 3792 12903 3844 12912
rect 3792 12869 3801 12903
rect 3801 12869 3835 12903
rect 3835 12869 3844 12903
rect 3792 12860 3844 12869
rect 5356 12928 5408 12980
rect 5540 12928 5592 12980
rect 6920 12928 6972 12980
rect 4988 12860 5040 12912
rect 6092 12860 6144 12912
rect 6828 12860 6880 12912
rect 9312 12928 9364 12980
rect 10600 12928 10652 12980
rect 1124 12792 1176 12844
rect 1492 12792 1544 12844
rect 3608 12792 3660 12844
rect 4068 12792 4120 12844
rect 2688 12724 2740 12776
rect 4160 12724 4212 12776
rect 6184 12792 6236 12844
rect 6736 12792 6788 12844
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6000 12724 6052 12733
rect 7748 12792 7800 12844
rect 10416 12860 10468 12912
rect 10508 12903 10560 12912
rect 10508 12869 10517 12903
rect 10517 12869 10551 12903
rect 10551 12869 10560 12903
rect 10508 12860 10560 12869
rect 10876 12860 10928 12912
rect 9496 12792 9548 12844
rect 10232 12792 10284 12844
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12716 12928 12768 12980
rect 15200 12928 15252 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17592 12971 17644 12980
rect 17592 12937 17601 12971
rect 17601 12937 17635 12971
rect 17635 12937 17644 12971
rect 17592 12928 17644 12937
rect 23296 12928 23348 12980
rect 13360 12792 13412 12844
rect 7656 12724 7708 12776
rect 6736 12656 6788 12708
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 7748 12588 7800 12640
rect 8392 12588 8444 12640
rect 10968 12588 11020 12640
rect 11336 12588 11388 12640
rect 12808 12724 12860 12776
rect 15476 12792 15528 12844
rect 12348 12656 12400 12708
rect 14924 12724 14976 12776
rect 18512 12792 18564 12844
rect 19524 12903 19576 12912
rect 19524 12869 19533 12903
rect 19533 12869 19567 12903
rect 19567 12869 19576 12903
rect 19524 12860 19576 12869
rect 20260 12903 20312 12912
rect 20260 12869 20269 12903
rect 20269 12869 20303 12903
rect 20303 12869 20312 12903
rect 20260 12860 20312 12869
rect 20720 12860 20772 12912
rect 22192 12860 22244 12912
rect 15936 12656 15988 12708
rect 12716 12588 12768 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 14372 12588 14424 12640
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 17040 12724 17092 12776
rect 17592 12724 17644 12776
rect 18236 12588 18288 12640
rect 18328 12631 18380 12640
rect 18328 12597 18337 12631
rect 18337 12597 18371 12631
rect 18371 12597 18380 12631
rect 18328 12588 18380 12597
rect 18972 12767 19024 12776
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 21088 12792 21140 12844
rect 21456 12792 21508 12844
rect 23204 12860 23256 12912
rect 23756 12860 23808 12912
rect 26240 12792 26292 12844
rect 26424 12724 26476 12776
rect 23388 12588 23440 12640
rect 24676 12588 24728 12640
rect 25872 12631 25924 12640
rect 25872 12597 25881 12631
rect 25881 12597 25915 12631
rect 25915 12597 25924 12631
rect 25872 12588 25924 12597
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2412 12384 2464 12436
rect 3608 12384 3660 12436
rect 4068 12384 4120 12436
rect 4896 12384 4948 12436
rect 7656 12384 7708 12436
rect 3424 12316 3476 12368
rect 3792 12248 3844 12300
rect 5448 12248 5500 12300
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 7196 12316 7248 12368
rect 10876 12384 10928 12436
rect 10968 12384 11020 12436
rect 14740 12384 14792 12436
rect 15384 12384 15436 12436
rect 18236 12384 18288 12436
rect 18788 12384 18840 12436
rect 6368 12248 6420 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3148 12180 3200 12232
rect 3240 12180 3292 12232
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 12072 12316 12124 12368
rect 9312 12248 9364 12300
rect 10876 12248 10928 12300
rect 14004 12316 14056 12368
rect 14096 12359 14148 12368
rect 14096 12325 14105 12359
rect 14105 12325 14139 12359
rect 14139 12325 14148 12359
rect 14096 12316 14148 12325
rect 17500 12316 17552 12368
rect 1952 12112 2004 12164
rect 8944 12180 8996 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 10232 12180 10284 12232
rect 4344 12044 4396 12096
rect 4988 12044 5040 12096
rect 6000 12044 6052 12096
rect 6552 12112 6604 12164
rect 7380 12112 7432 12164
rect 7472 12044 7524 12096
rect 7656 12112 7708 12164
rect 8392 12044 8444 12096
rect 10416 12112 10468 12164
rect 13820 12112 13872 12164
rect 14740 12180 14792 12232
rect 15200 12248 15252 12300
rect 17224 12248 17276 12300
rect 18328 12248 18380 12300
rect 16120 12180 16172 12232
rect 19064 12316 19116 12368
rect 22744 12384 22796 12436
rect 23296 12384 23348 12436
rect 25964 12384 26016 12436
rect 19524 12248 19576 12300
rect 22192 12248 22244 12300
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 23572 12316 23624 12368
rect 24952 12316 25004 12368
rect 24768 12248 24820 12300
rect 10784 12044 10836 12096
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 11888 12044 11940 12096
rect 12348 12044 12400 12096
rect 12440 12044 12492 12096
rect 12624 12044 12676 12096
rect 12808 12044 12860 12096
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 13912 12044 13964 12096
rect 14096 12044 14148 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 16488 12155 16540 12164
rect 16488 12121 16497 12155
rect 16497 12121 16531 12155
rect 16531 12121 16540 12155
rect 16488 12112 16540 12121
rect 17040 12112 17092 12164
rect 19432 12180 19484 12232
rect 19524 12112 19576 12164
rect 23664 12180 23716 12232
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 22560 12155 22612 12164
rect 22560 12121 22569 12155
rect 22569 12121 22603 12155
rect 22603 12121 22612 12155
rect 22560 12112 22612 12121
rect 24676 12112 24728 12164
rect 17868 12044 17920 12096
rect 20720 12044 20772 12096
rect 21364 12044 21416 12096
rect 21824 12087 21876 12096
rect 21824 12053 21833 12087
rect 21833 12053 21867 12087
rect 21867 12053 21876 12087
rect 21824 12044 21876 12053
rect 23848 12044 23900 12096
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 24400 12044 24452 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 2412 11840 2464 11892
rect 2872 11840 2924 11892
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 4712 11840 4764 11892
rect 5724 11840 5776 11892
rect 6000 11840 6052 11892
rect 7564 11840 7616 11892
rect 8024 11840 8076 11892
rect 10508 11840 10560 11892
rect 11888 11840 11940 11892
rect 13728 11840 13780 11892
rect 16304 11840 16356 11892
rect 7380 11772 7432 11824
rect 7932 11772 7984 11824
rect 9128 11772 9180 11824
rect 11060 11772 11112 11824
rect 2504 11704 2556 11756
rect 3884 11704 3936 11756
rect 5264 11704 5316 11756
rect 6552 11704 6604 11756
rect 5540 11636 5592 11688
rect 6092 11636 6144 11688
rect 6368 11636 6420 11688
rect 8944 11704 8996 11756
rect 13452 11815 13504 11824
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 14464 11772 14516 11824
rect 16856 11840 16908 11892
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 8392 11636 8444 11688
rect 12256 11636 12308 11688
rect 14740 11704 14792 11756
rect 16672 11704 16724 11756
rect 16948 11772 17000 11824
rect 17868 11704 17920 11756
rect 35348 11840 35400 11892
rect 20720 11772 20772 11824
rect 21364 11772 21416 11824
rect 21640 11772 21692 11824
rect 22284 11772 22336 11824
rect 22744 11772 22796 11824
rect 23664 11772 23716 11824
rect 25136 11704 25188 11756
rect 39304 11704 39356 11756
rect 3148 11568 3200 11620
rect 7196 11568 7248 11620
rect 8668 11568 8720 11620
rect 10692 11568 10744 11620
rect 1952 11500 2004 11552
rect 2872 11500 2924 11552
rect 3608 11500 3660 11552
rect 3884 11500 3936 11552
rect 6644 11500 6696 11552
rect 7472 11500 7524 11552
rect 12256 11500 12308 11552
rect 13820 11636 13872 11688
rect 16304 11636 16356 11688
rect 17040 11636 17092 11688
rect 17684 11636 17736 11688
rect 19524 11636 19576 11688
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 25872 11636 25924 11688
rect 13820 11500 13872 11552
rect 13912 11500 13964 11552
rect 15200 11500 15252 11552
rect 16396 11500 16448 11552
rect 18972 11500 19024 11552
rect 23940 11500 23992 11552
rect 24400 11543 24452 11552
rect 24400 11509 24409 11543
rect 24409 11509 24443 11543
rect 24443 11509 24452 11543
rect 24400 11500 24452 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 3700 11296 3752 11348
rect 3976 11296 4028 11348
rect 3608 11228 3660 11280
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 6920 11296 6972 11348
rect 7288 11296 7340 11348
rect 8668 11296 8720 11348
rect 7380 11228 7432 11280
rect 7932 11228 7984 11280
rect 8760 11228 8812 11280
rect 8024 11160 8076 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 2780 11092 2832 11144
rect 4896 11092 4948 11144
rect 7288 11092 7340 11144
rect 7840 11092 7892 11144
rect 9956 11228 10008 11280
rect 10416 11339 10468 11348
rect 10416 11305 10425 11339
rect 10425 11305 10459 11339
rect 10459 11305 10468 11339
rect 10416 11296 10468 11305
rect 12440 11296 12492 11348
rect 13360 11296 13412 11348
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 15660 11296 15712 11348
rect 16120 11296 16172 11348
rect 9312 11160 9364 11212
rect 11152 11160 11204 11212
rect 16396 11228 16448 11280
rect 19248 11296 19300 11348
rect 19984 11296 20036 11348
rect 18420 11228 18472 11280
rect 18972 11228 19024 11280
rect 22652 11271 22704 11280
rect 22652 11237 22661 11271
rect 22661 11237 22695 11271
rect 22695 11237 22704 11271
rect 22652 11228 22704 11237
rect 12256 11160 12308 11212
rect 13820 11160 13872 11212
rect 14648 11160 14700 11212
rect 16304 11160 16356 11212
rect 19248 11160 19300 11212
rect 25964 11160 26016 11212
rect 9680 11092 9732 11144
rect 9956 11092 10008 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12900 11092 12952 11144
rect 14372 11092 14424 11144
rect 17040 11092 17092 11144
rect 20628 11092 20680 11144
rect 24032 11092 24084 11144
rect 31300 11092 31352 11144
rect 5264 11067 5316 11076
rect 5264 11033 5273 11067
rect 5273 11033 5307 11067
rect 5307 11033 5316 11067
rect 5264 11024 5316 11033
rect 3608 10956 3660 11008
rect 5356 10956 5408 11008
rect 6276 10956 6328 11008
rect 7012 10956 7064 11008
rect 11796 11024 11848 11076
rect 11888 11067 11940 11076
rect 11888 11033 11897 11067
rect 11897 11033 11931 11067
rect 11931 11033 11940 11067
rect 11888 11024 11940 11033
rect 12624 11024 12676 11076
rect 15200 11024 15252 11076
rect 15568 11024 15620 11076
rect 17868 11024 17920 11076
rect 19432 11024 19484 11076
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 21640 11024 21692 11076
rect 23664 11024 23716 11076
rect 24400 11024 24452 11076
rect 27804 11024 27856 11076
rect 31392 11024 31444 11076
rect 47584 11092 47636 11144
rect 9772 10956 9824 11008
rect 13268 10956 13320 11008
rect 22100 10956 22152 11008
rect 24308 10956 24360 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1492 10795 1544 10804
rect 1492 10761 1501 10795
rect 1501 10761 1535 10795
rect 1535 10761 1544 10795
rect 1492 10752 1544 10761
rect 1860 10752 1912 10804
rect 3424 10795 3476 10804
rect 3424 10761 3433 10795
rect 3433 10761 3467 10795
rect 3467 10761 3476 10795
rect 3424 10752 3476 10761
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 5264 10752 5316 10804
rect 5908 10752 5960 10804
rect 6644 10752 6696 10804
rect 7196 10752 7248 10804
rect 2596 10684 2648 10736
rect 3516 10684 3568 10736
rect 480 10616 532 10668
rect 940 10616 992 10668
rect 1860 10616 1912 10668
rect 8300 10684 8352 10736
rect 8760 10684 8812 10736
rect 10968 10752 11020 10804
rect 11704 10752 11756 10804
rect 11980 10752 12032 10804
rect 12072 10752 12124 10804
rect 12348 10752 12400 10804
rect 13176 10752 13228 10804
rect 13268 10752 13320 10804
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 15752 10752 15804 10804
rect 10876 10684 10928 10736
rect 12716 10684 12768 10736
rect 12900 10684 12952 10736
rect 14464 10684 14516 10736
rect 17224 10684 17276 10736
rect 6276 10616 6328 10668
rect 5448 10548 5500 10600
rect 9588 10616 9640 10668
rect 5080 10480 5132 10532
rect 7380 10548 7432 10600
rect 6276 10412 6328 10464
rect 6644 10412 6696 10464
rect 8576 10548 8628 10600
rect 9036 10548 9088 10600
rect 11612 10616 11664 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 9128 10480 9180 10532
rect 10048 10480 10100 10532
rect 13728 10548 13780 10600
rect 11980 10480 12032 10532
rect 13544 10480 13596 10532
rect 16948 10616 17000 10668
rect 17132 10616 17184 10668
rect 19524 10752 19576 10804
rect 17868 10684 17920 10736
rect 21640 10752 21692 10804
rect 22560 10752 22612 10804
rect 16120 10548 16172 10600
rect 15936 10480 15988 10532
rect 8392 10412 8444 10464
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 12164 10412 12216 10464
rect 12624 10412 12676 10464
rect 12900 10412 12952 10464
rect 13176 10412 13228 10464
rect 16304 10548 16356 10600
rect 19064 10548 19116 10600
rect 18880 10480 18932 10532
rect 21272 10684 21324 10736
rect 21824 10616 21876 10668
rect 22652 10616 22704 10668
rect 18420 10412 18472 10464
rect 19524 10412 19576 10464
rect 20628 10412 20680 10464
rect 24308 10412 24360 10464
rect 34888 10412 34940 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 388 10208 440 10260
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 4068 10208 4120 10260
rect 4528 10208 4580 10260
rect 6552 10208 6604 10260
rect 13544 10208 13596 10260
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 17224 10208 17276 10260
rect 20168 10208 20220 10260
rect 22192 10208 22244 10260
rect 1400 10072 1452 10124
rect 1032 10004 1084 10056
rect 296 9868 348 9920
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 5264 9936 5316 9988
rect 7472 10140 7524 10192
rect 6000 10072 6052 10124
rect 7748 10072 7800 10124
rect 14372 10140 14424 10192
rect 16396 10183 16448 10192
rect 16396 10149 16405 10183
rect 16405 10149 16439 10183
rect 16439 10149 16448 10183
rect 16396 10140 16448 10149
rect 9864 10072 9916 10124
rect 14648 10115 14700 10124
rect 14648 10081 14657 10115
rect 14657 10081 14691 10115
rect 14691 10081 14700 10115
rect 14648 10072 14700 10081
rect 14924 10072 14976 10124
rect 16304 10072 16356 10124
rect 16856 10072 16908 10124
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 19524 10115 19576 10124
rect 19524 10081 19533 10115
rect 19533 10081 19567 10115
rect 19567 10081 19576 10115
rect 19524 10072 19576 10081
rect 22652 10072 22704 10124
rect 8392 9936 8444 9988
rect 9404 9979 9456 9988
rect 9404 9945 9413 9979
rect 9413 9945 9447 9979
rect 9447 9945 9456 9979
rect 9404 9936 9456 9945
rect 9864 9936 9916 9988
rect 21272 10004 21324 10056
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 24676 10004 24728 10056
rect 11612 9936 11664 9988
rect 11796 9936 11848 9988
rect 6920 9868 6972 9920
rect 7748 9868 7800 9920
rect 10324 9868 10376 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 11152 9868 11204 9920
rect 11980 9868 12032 9920
rect 12164 9936 12216 9988
rect 15200 9936 15252 9988
rect 12716 9868 12768 9920
rect 13268 9868 13320 9920
rect 13636 9868 13688 9920
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 15568 9868 15620 9920
rect 17868 9936 17920 9988
rect 18696 9868 18748 9920
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 1676 9596 1728 9648
rect 2136 9596 2188 9648
rect 3332 9639 3384 9648
rect 3332 9605 3341 9639
rect 3341 9605 3375 9639
rect 3375 9605 3384 9639
rect 3332 9596 3384 9605
rect 4252 9596 4304 9648
rect 5080 9596 5132 9648
rect 6000 9639 6052 9648
rect 6000 9605 6009 9639
rect 6009 9605 6043 9639
rect 6043 9605 6052 9639
rect 6000 9596 6052 9605
rect 2596 9392 2648 9444
rect 3424 9528 3476 9580
rect 3884 9528 3936 9580
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 5172 9528 5224 9580
rect 5448 9528 5500 9580
rect 7012 9596 7064 9648
rect 9312 9664 9364 9716
rect 10508 9664 10560 9716
rect 10876 9664 10928 9716
rect 8760 9596 8812 9648
rect 8944 9596 8996 9648
rect 10692 9639 10744 9648
rect 10692 9605 10701 9639
rect 10701 9605 10735 9639
rect 10735 9605 10744 9639
rect 10692 9596 10744 9605
rect 11152 9664 11204 9716
rect 14280 9664 14332 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 22744 9664 22796 9716
rect 24584 9664 24636 9716
rect 11980 9596 12032 9648
rect 13636 9596 13688 9648
rect 11612 9528 11664 9580
rect 13268 9528 13320 9580
rect 15108 9596 15160 9648
rect 15568 9596 15620 9648
rect 17224 9596 17276 9648
rect 18696 9596 18748 9648
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 18512 9528 18564 9580
rect 3424 9435 3476 9444
rect 3424 9401 3433 9435
rect 3433 9401 3467 9435
rect 3467 9401 3476 9435
rect 3424 9392 3476 9401
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 8300 9460 8352 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 6920 9324 6972 9376
rect 9864 9460 9916 9512
rect 11152 9460 11204 9512
rect 11980 9503 12032 9512
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 12348 9460 12400 9512
rect 14188 9460 14240 9512
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 15384 9460 15436 9512
rect 10048 9324 10100 9376
rect 11704 9392 11756 9444
rect 10876 9324 10928 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 17316 9324 17368 9376
rect 18972 9460 19024 9512
rect 20904 9639 20956 9648
rect 20904 9605 20913 9639
rect 20913 9605 20947 9639
rect 20947 9605 20956 9639
rect 20904 9596 20956 9605
rect 22100 9596 22152 9648
rect 22652 9639 22704 9648
rect 22652 9605 22661 9639
rect 22661 9605 22695 9639
rect 22695 9605 22704 9639
rect 22652 9596 22704 9605
rect 27804 9639 27856 9648
rect 27804 9605 27813 9639
rect 27813 9605 27847 9639
rect 27847 9605 27856 9639
rect 27804 9596 27856 9605
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 23940 9528 23992 9580
rect 24032 9528 24084 9580
rect 21272 9460 21324 9512
rect 26056 9392 26108 9444
rect 19156 9324 19208 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 1400 9120 1452 9172
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 4712 9163 4764 9172
rect 4712 9129 4721 9163
rect 4721 9129 4755 9163
rect 4755 9129 4764 9163
rect 4712 9120 4764 9129
rect 4896 9120 4948 9172
rect 1676 9052 1728 9104
rect 2504 9052 2556 9104
rect 6184 9120 6236 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 7656 9120 7708 9172
rect 10140 9120 10192 9172
rect 1216 8984 1268 9036
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 7472 9052 7524 9104
rect 3976 8916 4028 8968
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 5356 8916 5408 8968
rect 7104 8984 7156 9036
rect 7840 8984 7892 9036
rect 8760 9052 8812 9104
rect 9588 9052 9640 9104
rect 13360 9120 13412 9172
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7656 8916 7708 8968
rect 8668 8916 8720 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10324 8984 10376 9036
rect 10140 8916 10192 8968
rect 10692 8916 10744 8968
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 11704 8984 11756 9036
rect 12808 8984 12860 9036
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13360 8984 13412 9036
rect 13912 8984 13964 9036
rect 12716 8916 12768 8968
rect 4252 8891 4304 8900
rect 4252 8857 4261 8891
rect 4261 8857 4295 8891
rect 4295 8857 4304 8891
rect 4252 8848 4304 8857
rect 4344 8848 4396 8900
rect 8484 8848 8536 8900
rect 2504 8780 2556 8832
rect 2688 8780 2740 8832
rect 5172 8780 5224 8832
rect 7380 8780 7432 8832
rect 9588 8848 9640 8900
rect 9864 8848 9916 8900
rect 12164 8848 12216 8900
rect 12256 8848 12308 8900
rect 14188 8848 14240 8900
rect 15568 9052 15620 9104
rect 17776 9120 17828 9172
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 21180 9120 21232 9172
rect 31392 9120 31444 9172
rect 21732 9052 21784 9104
rect 16856 8984 16908 9036
rect 24768 8984 24820 9036
rect 35440 8984 35492 9036
rect 18328 8916 18380 8968
rect 21272 8916 21324 8968
rect 9036 8780 9088 8832
rect 10876 8780 10928 8832
rect 11336 8780 11388 8832
rect 11796 8780 11848 8832
rect 12532 8780 12584 8832
rect 13636 8780 13688 8832
rect 15108 8780 15160 8832
rect 16580 8848 16632 8900
rect 16764 8848 16816 8900
rect 20536 8848 20588 8900
rect 17776 8823 17828 8832
rect 17776 8789 17785 8823
rect 17785 8789 17819 8823
rect 17819 8789 17828 8823
rect 17776 8780 17828 8789
rect 19524 8823 19576 8832
rect 19524 8789 19533 8823
rect 19533 8789 19567 8823
rect 19567 8789 19576 8823
rect 19524 8780 19576 8789
rect 26240 8780 26292 8832
rect 28724 8780 28776 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 1768 8576 1820 8628
rect 1860 8440 1912 8492
rect 4804 8576 4856 8628
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5908 8576 5960 8628
rect 6184 8576 6236 8628
rect 9680 8576 9732 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 10416 8576 10468 8628
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 12808 8576 12860 8628
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 16488 8576 16540 8628
rect 16580 8576 16632 8628
rect 18696 8576 18748 8628
rect 19248 8619 19300 8628
rect 19248 8585 19257 8619
rect 19257 8585 19291 8619
rect 19291 8585 19300 8619
rect 19248 8576 19300 8585
rect 2044 8508 2096 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 4344 8508 4396 8560
rect 4620 8508 4672 8560
rect 6000 8508 6052 8560
rect 6276 8508 6328 8560
rect 3424 8440 3476 8492
rect 4988 8440 5040 8492
rect 2136 8372 2188 8424
rect 5448 8372 5500 8424
rect 6736 8440 6788 8492
rect 7564 8440 7616 8492
rect 9404 8551 9456 8560
rect 9404 8517 9413 8551
rect 9413 8517 9447 8551
rect 9447 8517 9456 8551
rect 9404 8508 9456 8517
rect 9588 8508 9640 8560
rect 10508 8508 10560 8560
rect 8668 8440 8720 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 7656 8372 7708 8424
rect 7840 8372 7892 8424
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 3148 8304 3200 8356
rect 6644 8304 6696 8356
rect 7564 8304 7616 8356
rect 9864 8372 9916 8424
rect 11428 8508 11480 8560
rect 12532 8508 12584 8560
rect 14188 8440 14240 8492
rect 14280 8440 14332 8492
rect 22008 8508 22060 8560
rect 8300 8304 8352 8356
rect 11060 8304 11112 8356
rect 11612 8304 11664 8356
rect 12348 8304 12400 8356
rect 6276 8236 6328 8288
rect 7840 8236 7892 8288
rect 12716 8236 12768 8288
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 16120 8440 16172 8492
rect 17316 8440 17368 8492
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 15568 8372 15620 8424
rect 16764 8372 16816 8424
rect 16856 8372 16908 8424
rect 17592 8440 17644 8492
rect 18880 8440 18932 8492
rect 18696 8372 18748 8424
rect 19432 8372 19484 8424
rect 13912 8304 13964 8356
rect 19524 8347 19576 8356
rect 19524 8313 19533 8347
rect 19533 8313 19567 8347
rect 19567 8313 19576 8347
rect 19524 8304 19576 8313
rect 16856 8236 16908 8288
rect 23664 8236 23716 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 2136 8032 2188 8084
rect 2504 8032 2556 8084
rect 7012 8032 7064 8084
rect 7564 8032 7616 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 9680 8032 9732 8084
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 13636 8032 13688 8084
rect 14740 8032 14792 8084
rect 14832 8032 14884 8084
rect 17408 8032 17460 8084
rect 756 7964 808 8016
rect 2412 7896 2464 7948
rect 1308 7828 1360 7880
rect 7656 7964 7708 8016
rect 5724 7896 5776 7948
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5540 7828 5592 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 9864 7964 9916 8016
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 3240 7692 3292 7744
rect 6736 7760 6788 7812
rect 7472 7760 7524 7812
rect 9864 7828 9916 7880
rect 11336 7964 11388 8016
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 10692 7828 10744 7880
rect 11244 7828 11296 7880
rect 12440 7760 12492 7812
rect 12716 7896 12768 7948
rect 17132 7896 17184 7948
rect 13452 7828 13504 7880
rect 14188 7828 14240 7880
rect 16028 7828 16080 7880
rect 15292 7760 15344 7812
rect 16212 7828 16264 7880
rect 18420 7828 18472 7880
rect 17776 7760 17828 7812
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 6920 7692 6972 7744
rect 7380 7692 7432 7744
rect 8668 7692 8720 7744
rect 10048 7692 10100 7744
rect 11060 7692 11112 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 5356 7488 5408 7540
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 6276 7488 6328 7540
rect 10784 7488 10836 7540
rect 11060 7488 11112 7540
rect 12072 7488 12124 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 15200 7488 15252 7540
rect 24032 7531 24084 7540
rect 24032 7497 24041 7531
rect 24041 7497 24075 7531
rect 24075 7497 24084 7531
rect 24032 7488 24084 7497
rect 2228 7352 2280 7404
rect 6276 7352 6328 7404
rect 7104 7352 7156 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7472 7352 7524 7404
rect 7840 7352 7892 7404
rect 8668 7352 8720 7404
rect 8944 7352 8996 7404
rect 10508 7352 10560 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 12348 7352 12400 7404
rect 13360 7352 13412 7404
rect 13820 7352 13872 7404
rect 2872 7327 2924 7336
rect 2872 7293 2881 7327
rect 2881 7293 2915 7327
rect 2915 7293 2924 7327
rect 2872 7284 2924 7293
rect 4712 7284 4764 7336
rect 5632 7284 5684 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 6920 7284 6972 7336
rect 8760 7284 8812 7336
rect 664 7148 716 7200
rect 6184 7216 6236 7268
rect 7012 7148 7064 7200
rect 10232 7259 10284 7268
rect 10232 7225 10241 7259
rect 10241 7225 10275 7259
rect 10275 7225 10284 7259
rect 10232 7216 10284 7225
rect 11520 7284 11572 7336
rect 15108 7420 15160 7472
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 20628 7352 20680 7404
rect 23664 7352 23716 7404
rect 21088 7284 21140 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 16028 7216 16080 7268
rect 7840 7148 7892 7200
rect 12164 7148 12216 7200
rect 12348 7191 12400 7200
rect 12348 7157 12357 7191
rect 12357 7157 12391 7191
rect 12391 7157 12400 7191
rect 12348 7148 12400 7157
rect 13360 7148 13412 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 112 6876 164 6928
rect 6828 6944 6880 6996
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 7380 6944 7432 6996
rect 7840 6944 7892 6996
rect 5632 6876 5684 6928
rect 15936 6876 15988 6928
rect 1952 6808 2004 6860
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 3240 6808 3292 6860
rect 2780 6740 2832 6792
rect 3700 6740 3752 6792
rect 4160 6808 4212 6860
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 1308 6672 1360 6724
rect 480 6604 532 6656
rect 5080 6672 5132 6724
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 11888 6808 11940 6860
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 7840 6740 7892 6792
rect 5540 6604 5592 6656
rect 6920 6604 6972 6656
rect 7104 6604 7156 6656
rect 8484 6672 8536 6724
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 11612 6740 11664 6792
rect 11796 6740 11848 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 22560 6808 22612 6860
rect 20720 6783 20772 6792
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 10508 6715 10560 6724
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 10876 6715 10928 6724
rect 10876 6681 10885 6715
rect 10885 6681 10919 6715
rect 10919 6681 10928 6715
rect 10876 6672 10928 6681
rect 10784 6604 10836 6656
rect 12348 6672 12400 6724
rect 14096 6604 14148 6656
rect 18512 6604 18564 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 1308 6264 1360 6316
rect 3240 6332 3292 6384
rect 3608 6400 3660 6452
rect 4068 6400 4120 6452
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 6000 6400 6052 6452
rect 6828 6400 6880 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 10600 6400 10652 6452
rect 11428 6400 11480 6452
rect 14648 6400 14700 6452
rect 5356 6332 5408 6384
rect 21916 6332 21968 6384
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 4344 6264 4396 6316
rect 572 6196 624 6248
rect 9404 6264 9456 6316
rect 9496 6264 9548 6316
rect 10416 6264 10468 6316
rect 11704 6264 11756 6316
rect 12348 6264 12400 6316
rect 12808 6264 12860 6316
rect 22284 6264 22336 6316
rect 28724 6332 28776 6384
rect 6644 6196 6696 6248
rect 9680 6196 9732 6248
rect 11980 6196 12032 6248
rect 4436 6128 4488 6180
rect 7012 6128 7064 6180
rect 14004 6128 14056 6180
rect 1860 6060 1912 6112
rect 4160 6060 4212 6112
rect 6920 6060 6972 6112
rect 7104 6060 7156 6112
rect 16672 6060 16724 6112
rect 24032 6128 24084 6180
rect 23572 6060 23624 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 2504 5856 2556 5908
rect 9036 5856 9088 5908
rect 9312 5856 9364 5908
rect 9772 5856 9824 5908
rect 16856 5856 16908 5908
rect 19524 5856 19576 5908
rect 6368 5788 6420 5840
rect 7748 5788 7800 5840
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 3516 5720 3568 5772
rect 3976 5720 4028 5772
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 3516 5584 3568 5636
rect 3884 5584 3936 5636
rect 2320 5516 2372 5568
rect 4620 5652 4672 5704
rect 6552 5720 6604 5772
rect 9128 5652 9180 5704
rect 13728 5720 13780 5772
rect 14556 5720 14608 5772
rect 14740 5720 14792 5772
rect 17040 5720 17092 5772
rect 20720 5720 20772 5772
rect 6736 5584 6788 5636
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 6460 5516 6512 5568
rect 10692 5516 10744 5568
rect 15108 5516 15160 5568
rect 16304 5584 16356 5636
rect 19432 5584 19484 5636
rect 26240 5856 26292 5908
rect 23480 5720 23532 5772
rect 26700 5763 26752 5772
rect 26700 5729 26709 5763
rect 26709 5729 26743 5763
rect 26743 5729 26752 5763
rect 26700 5720 26752 5729
rect 24768 5584 24820 5636
rect 27528 5584 27580 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 4068 5312 4120 5364
rect 5724 5312 5776 5364
rect 3792 5244 3844 5296
rect 4436 5244 4488 5296
rect 4528 5176 4580 5228
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 22284 5312 22336 5364
rect 23480 5312 23532 5364
rect 24768 5244 24820 5296
rect 27620 5244 27672 5296
rect 28540 5244 28592 5296
rect 29092 5244 29144 5296
rect 20904 5176 20956 5185
rect 23572 5176 23624 5228
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 6092 5040 6144 5092
rect 18604 5040 18656 5092
rect 21364 5083 21416 5092
rect 21364 5049 21373 5083
rect 21373 5049 21407 5083
rect 21407 5049 21416 5083
rect 21364 5040 21416 5049
rect 25504 5040 25556 5092
rect 27344 5151 27396 5160
rect 27344 5117 27353 5151
rect 27353 5117 27387 5151
rect 27387 5117 27396 5151
rect 27344 5108 27396 5117
rect 29092 5040 29144 5092
rect 29644 5151 29696 5160
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 31760 5108 31812 5160
rect 32496 5108 32548 5160
rect 32864 5040 32916 5092
rect 4988 4972 5040 5024
rect 20720 4972 20772 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 3332 4768 3384 4820
rect 3516 4768 3568 4820
rect 3792 4768 3844 4820
rect 4068 4768 4120 4820
rect 10140 4768 10192 4820
rect 16304 4768 16356 4820
rect 9956 4700 10008 4752
rect 27344 4768 27396 4820
rect 1308 4632 1360 4684
rect 4712 4632 4764 4684
rect 2596 4564 2648 4616
rect 3424 4564 3476 4616
rect 4252 4564 4304 4616
rect 11060 4564 11112 4616
rect 29644 4700 29696 4752
rect 15108 4632 15160 4684
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 19892 4632 19944 4684
rect 20904 4564 20956 4616
rect 21364 4564 21416 4616
rect 8852 4496 8904 4548
rect 13820 4496 13872 4548
rect 23572 4496 23624 4548
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 2044 4088 2096 4140
rect 2780 4088 2832 4140
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 14096 4020 14148 4072
rect 18604 4020 18656 4072
rect 20076 4020 20128 4072
rect 388 3952 440 4004
rect 8944 3952 8996 4004
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 2780 3680 2832 3732
rect 7564 3680 7616 3732
rect 12440 3680 12492 3732
rect 13728 3680 13780 3732
rect 32496 3680 32548 3732
rect 41420 3680 41472 3732
rect 2872 3655 2924 3664
rect 2872 3621 2881 3655
rect 2881 3621 2915 3655
rect 2915 3621 2924 3655
rect 2872 3612 2924 3621
rect 3424 3655 3476 3664
rect 3424 3621 3433 3655
rect 3433 3621 3467 3655
rect 3467 3621 3476 3655
rect 3424 3612 3476 3621
rect 29184 3612 29236 3664
rect 44088 3612 44140 3664
rect 1308 3544 1360 3596
rect 26700 3544 26752 3596
rect 46756 3544 46808 3596
rect 3332 3476 3384 3528
rect 4068 3476 4120 3528
rect 27620 3476 27672 3528
rect 49424 3476 49476 3528
rect 7472 3408 7524 3460
rect 19340 3408 19392 3460
rect 38752 3408 38804 3460
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 3240 3136 3292 3188
rect 1216 3068 1268 3120
rect 8300 3136 8352 3188
rect 2872 3000 2924 3052
rect 8760 3068 8812 3120
rect 11060 3136 11112 3188
rect 12440 3068 12492 3120
rect 13820 3068 13872 3120
rect 14096 3111 14148 3120
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 19892 3068 19944 3120
rect 8392 3000 8444 3052
rect 10140 3000 10192 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 1308 2864 1360 2916
rect 7380 2932 7432 2984
rect 8024 2932 8076 2984
rect 9772 2932 9824 2984
rect 22744 2932 22796 2984
rect 1400 2796 1452 2848
rect 2780 2796 2832 2848
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 12440 2796 12492 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 1308 2456 1360 2508
rect 4344 2592 4396 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27528 2592 27580 2644
rect 29092 2592 29144 2644
rect 32864 2592 32916 2644
rect 15016 2524 15068 2576
rect 1216 2388 1268 2440
rect 2872 2456 2924 2508
rect 4068 2456 4120 2508
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 12072 2456 12124 2508
rect 28724 2456 28776 2508
rect 2780 2388 2832 2440
rect 8300 2388 8352 2440
rect 9772 2388 9824 2440
rect 12440 2388 12492 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 11888 2320 11940 2372
rect 8024 2252 8076 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 1308 2048 1360 2100
rect 3332 2048 3384 2100
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26330 2926 27000
rect 2870 26302 3464 26330
rect 2870 26200 2926 26302
rect 1584 24336 1636 24342
rect 1582 24304 1584 24313
rect 1636 24304 1638 24313
rect 1582 24239 1638 24248
rect 1768 24200 1820 24206
rect 1766 24168 1768 24177
rect 2136 24200 2188 24206
rect 1820 24168 1822 24177
rect 756 24132 808 24138
rect 2136 24142 2188 24148
rect 1766 24103 1822 24112
rect 756 24074 808 24080
rect 572 23520 624 23526
rect 572 23462 624 23468
rect 480 20800 532 20806
rect 480 20742 532 20748
rect 492 16574 520 20742
rect 308 16546 520 16574
rect 204 15156 256 15162
rect 204 15098 256 15104
rect 112 13932 164 13938
rect 112 13874 164 13880
rect 124 6934 152 13874
rect 112 6928 164 6934
rect 216 6914 244 15098
rect 308 9926 336 16546
rect 584 16402 612 23462
rect 664 22772 716 22778
rect 664 22714 716 22720
rect 400 16374 612 16402
rect 400 10266 428 16374
rect 480 16244 532 16250
rect 480 16186 532 16192
rect 492 11642 520 16186
rect 492 11614 612 11642
rect 480 10668 532 10674
rect 480 10610 532 10616
rect 388 10260 440 10266
rect 388 10202 440 10208
rect 296 9920 348 9926
rect 296 9862 348 9868
rect 216 6886 428 6914
rect 112 6870 164 6876
rect 400 4010 428 6886
rect 492 6662 520 10610
rect 480 6656 532 6662
rect 480 6598 532 6604
rect 584 6254 612 11614
rect 676 7206 704 22714
rect 768 13938 796 24074
rect 848 23656 900 23662
rect 848 23598 900 23604
rect 756 13932 808 13938
rect 756 13874 808 13880
rect 756 13796 808 13802
rect 756 13738 808 13744
rect 768 8022 796 13738
rect 860 13410 888 23598
rect 940 22976 992 22982
rect 940 22918 992 22924
rect 952 13546 980 22918
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1124 21412 1176 21418
rect 1124 21354 1176 21360
rect 1032 20596 1084 20602
rect 1032 20538 1084 20544
rect 1044 13682 1072 20538
rect 1136 16946 1164 21354
rect 1320 20777 1348 22034
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1858 20496 1914 20505
rect 1858 20431 1914 20440
rect 1952 20460 2004 20466
rect 1674 19680 1730 19689
rect 1674 19615 1730 19624
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17921 1440 18770
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 1400 17604 1452 17610
rect 1400 17546 1452 17552
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1136 16918 1256 16946
rect 1122 16416 1178 16425
rect 1122 16351 1178 16360
rect 1136 16250 1164 16351
rect 1124 16244 1176 16250
rect 1124 16186 1176 16192
rect 1122 16144 1178 16153
rect 1122 16079 1178 16088
rect 1136 15162 1164 16079
rect 1124 15156 1176 15162
rect 1124 15098 1176 15104
rect 1122 15056 1178 15065
rect 1122 14991 1178 15000
rect 1136 14958 1164 14991
rect 1124 14952 1176 14958
rect 1124 14894 1176 14900
rect 1228 13802 1256 16918
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1216 13796 1268 13802
rect 1216 13738 1268 13744
rect 1044 13654 1348 13682
rect 952 13518 1256 13546
rect 1122 13424 1178 13433
rect 860 13382 1072 13410
rect 938 10704 994 10713
rect 938 10639 940 10648
rect 992 10639 994 10648
rect 940 10610 992 10616
rect 1044 10062 1072 13382
rect 1122 13359 1178 13368
rect 1136 12850 1164 13359
rect 1124 12844 1176 12850
rect 1124 12786 1176 12792
rect 1032 10056 1084 10062
rect 1032 9998 1084 10004
rect 1228 9042 1256 13518
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 756 8016 808 8022
rect 756 7958 808 7964
rect 1320 7886 1348 13654
rect 1412 10130 1440 17546
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 10810 1532 12786
rect 1688 12238 1716 19615
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1780 17202 1808 19450
rect 1872 18766 1900 20431
rect 1952 20402 2004 20408
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1766 13424 1822 13433
rect 1766 13359 1822 13368
rect 1780 13326 1808 13359
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1766 12200 1822 12209
rect 1584 11144 1636 11150
rect 1582 11112 1584 11121
rect 1636 11112 1638 11121
rect 1582 11047 1638 11056
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 9178 1440 10066
rect 1688 9654 1716 12174
rect 1964 12170 1992 20402
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2056 17513 2084 18158
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 2056 13394 2084 13767
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1766 12135 1822 12144
rect 1952 12164 2004 12170
rect 1492 9648 1544 9654
rect 1490 9616 1492 9625
rect 1676 9648 1728 9654
rect 1544 9616 1546 9625
rect 1676 9590 1728 9596
rect 1490 9551 1546 9560
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1688 9110 1716 9318
rect 1676 9104 1728 9110
rect 1676 9046 1728 9052
rect 1780 8974 1808 12135
rect 1952 12106 2004 12112
rect 1858 11656 1914 11665
rect 1858 11591 1914 11600
rect 1872 11218 1900 11591
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1872 10810 1900 10911
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1858 10704 1914 10713
rect 1858 10639 1860 10648
rect 1912 10639 1914 10648
rect 1860 10610 1912 10616
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1780 8634 1808 8910
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1872 8498 1900 10610
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 664 7200 716 7206
rect 664 7142 716 7148
rect 1964 6866 1992 11494
rect 2042 11112 2098 11121
rect 2042 11047 2098 11056
rect 2056 9178 2084 11047
rect 2148 9654 2176 24142
rect 2240 18426 2268 26200
rect 3146 25256 3202 25265
rect 3146 25191 3202 25200
rect 3160 24886 3188 25191
rect 3148 24880 3200 24886
rect 3148 24822 3200 24828
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2778 24440 2834 24449
rect 2950 24443 3258 24452
rect 2778 24375 2834 24384
rect 2792 24342 2820 24375
rect 2780 24336 2832 24342
rect 2780 24278 2832 24284
rect 3436 24154 3464 26302
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5304 26330
rect 4802 26200 4858 26302
rect 3528 24274 3556 26200
rect 3882 25664 3938 25673
rect 3882 25599 3938 25608
rect 3896 25226 3924 25599
rect 3884 25220 3936 25226
rect 3884 25162 3936 25168
rect 3698 24848 3754 24857
rect 3698 24783 3754 24792
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3436 24126 3648 24154
rect 2412 23792 2464 23798
rect 2412 23734 2464 23740
rect 2424 23526 2452 23734
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 3514 22536 3570 22545
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2320 21548 2372 21554
rect 2686 21519 2742 21528
rect 2320 21490 2372 21496
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6322 1348 6666
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 572 6248 624 6254
rect 572 6190 624 6196
rect 1320 6089 1348 6258
rect 1860 6112 1912 6118
rect 1306 6080 1362 6089
rect 1860 6054 1912 6060
rect 1306 6015 1362 6024
rect 1872 5778 1900 6054
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1320 4690 1348 5199
rect 1596 5166 1624 5607
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1582 4856 1638 4865
rect 1582 4791 1638 4800
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1596 4146 1624 4791
rect 2056 4146 2084 8502
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 8090 2176 8366
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2240 7410 2268 16594
rect 2332 8498 2360 21490
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 3514 22471 3570 22480
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3240 21616 3292 21622
rect 3436 21593 3464 21830
rect 3240 21558 3292 21564
rect 3422 21584 3478 21593
rect 3252 21350 3280 21558
rect 3422 21519 3478 21528
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2424 12442 2452 20266
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2516 12345 2544 19790
rect 2792 19530 2820 20334
rect 2884 19904 2912 20810
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19961 3372 21422
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3330 19952 3386 19961
rect 2884 19876 3004 19904
rect 3330 19887 3386 19896
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2700 19502 2820 19530
rect 2700 19145 2728 19502
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2686 19136 2742 19145
rect 2686 19071 2742 19080
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2502 12336 2558 12345
rect 2502 12271 2558 12280
rect 2410 11928 2466 11937
rect 2410 11863 2412 11872
rect 2464 11863 2466 11872
rect 2412 11834 2464 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2410 10432 2466 10441
rect 2410 10367 2466 10376
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2318 8120 2374 8129
rect 2318 8055 2374 8064
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2332 5574 2360 8055
rect 2424 7954 2452 10367
rect 2516 9110 2544 11698
rect 2608 10742 2636 18799
rect 2792 18329 2820 19314
rect 2884 18737 2912 19722
rect 2976 19553 3004 19876
rect 2962 19544 3018 19553
rect 2962 19479 3018 19488
rect 3330 19272 3386 19281
rect 3330 19207 3332 19216
rect 3384 19207 3386 19216
rect 3332 19178 3384 19184
rect 3436 19122 3464 21286
rect 3528 21010 3556 22471
rect 3620 21486 3648 24126
rect 3712 23662 3740 24783
rect 3974 24712 4030 24721
rect 3974 24647 4030 24656
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 3700 23656 3752 23662
rect 3700 23598 3752 23604
rect 3804 22386 3832 24550
rect 3988 24410 4016 24647
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3976 24132 4028 24138
rect 3976 24074 4028 24080
rect 3988 23633 4016 24074
rect 4066 24032 4122 24041
rect 4066 23967 4122 23976
rect 3974 23624 4030 23633
rect 4080 23610 4108 23967
rect 4172 23730 4200 26200
rect 4436 24880 4488 24886
rect 4250 24848 4306 24857
rect 4436 24822 4488 24828
rect 4250 24783 4306 24792
rect 4264 24410 4292 24783
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4356 24410 4384 24686
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4080 23582 4292 23610
rect 3974 23559 4030 23568
rect 3882 23216 3938 23225
rect 3882 23151 3938 23160
rect 3896 22522 3924 23151
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 4066 23080 4122 23089
rect 3988 22681 4016 23054
rect 4066 23015 4122 23024
rect 4080 22930 4108 23015
rect 4080 22902 4200 22930
rect 4066 22808 4122 22817
rect 4066 22743 4122 22752
rect 3974 22672 4030 22681
rect 3974 22607 4030 22616
rect 3896 22494 4016 22522
rect 3804 22358 3924 22386
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3712 22001 3740 22034
rect 3698 21992 3754 22001
rect 3698 21927 3754 21936
rect 3804 21729 3832 22102
rect 3790 21720 3846 21729
rect 3790 21655 3846 21664
rect 3700 21616 3752 21622
rect 3700 21558 3752 21564
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3516 21004 3568 21010
rect 3516 20946 3568 20952
rect 3606 20904 3662 20913
rect 3606 20839 3662 20848
rect 3620 20806 3648 20839
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3712 20482 3740 21558
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3344 19094 3464 19122
rect 3528 20454 3740 20482
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2870 18728 2926 18737
rect 2870 18663 2926 18672
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3344 17785 3372 19094
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3436 17882 3464 18906
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3330 17776 3386 17785
rect 3330 17711 3386 17720
rect 3528 17354 3556 20454
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3606 20224 3662 20233
rect 3606 20159 3662 20168
rect 3620 20058 3648 20159
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3712 19446 3740 20266
rect 3804 20244 3832 21082
rect 3896 21026 3924 22358
rect 3988 21146 4016 22494
rect 4080 22234 4108 22743
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4172 22114 4200 22902
rect 4080 22086 4200 22114
rect 4080 22030 4108 22086
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4172 21690 4200 21898
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 3896 20998 4108 21026
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 3936 20360 3938 20369
rect 3882 20295 3938 20304
rect 3804 20216 3924 20244
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3700 19440 3752 19446
rect 3606 19408 3662 19417
rect 3700 19382 3752 19388
rect 3606 19343 3608 19352
rect 3660 19343 3662 19352
rect 3608 19314 3660 19320
rect 3804 19258 3832 19450
rect 3712 19230 3832 19258
rect 3606 19136 3662 19145
rect 3606 19071 3662 19080
rect 3620 18902 3648 19071
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 2792 17326 3556 17354
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 12782 2728 15302
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2792 11506 2820 17326
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 11898 2912 17070
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3436 16697 3464 16730
rect 3422 16688 3478 16697
rect 3332 16652 3384 16658
rect 3422 16623 3478 16632
rect 3332 16594 3384 16600
rect 3344 16114 3372 16594
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 3516 15496 3568 15502
rect 3422 15464 3478 15473
rect 3516 15438 3568 15444
rect 3422 15399 3478 15408
rect 3436 15026 3464 15399
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3238 13016 3294 13025
rect 3344 12986 3372 14214
rect 3528 14074 3556 15438
rect 3606 14512 3662 14521
rect 3606 14447 3608 14456
rect 3660 14447 3662 14456
rect 3608 14418 3660 14424
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3514 13968 3570 13977
rect 3514 13903 3570 13912
rect 3608 13932 3660 13938
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3238 12951 3294 12960
rect 3332 12980 3384 12986
rect 3252 12866 3280 12951
rect 3332 12922 3384 12928
rect 3252 12838 3372 12866
rect 3344 12617 3372 12838
rect 3330 12608 3386 12617
rect 2950 12540 3258 12549
rect 3330 12543 3386 12552
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3436 12434 3464 13398
rect 3344 12406 3464 12434
rect 3148 12232 3200 12238
rect 3240 12232 3292 12238
rect 3148 12174 3200 12180
rect 3238 12200 3240 12209
rect 3292 12200 3294 12209
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2884 11558 2912 11834
rect 3160 11626 3188 12174
rect 3238 12135 3294 12144
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 2700 11478 2820 11506
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2700 11234 2728 11478
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2700 11206 2820 11234
rect 2792 11150 2820 11206
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2792 9674 2820 11086
rect 2870 10840 2926 10849
rect 2870 10775 2926 10784
rect 2700 9646 2820 9674
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8090 2544 8774
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2516 5914 2544 8026
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2608 4622 2636 9386
rect 2700 8838 2728 9646
rect 2778 9344 2834 9353
rect 2778 9279 2834 9288
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2792 7936 2820 9279
rect 2700 7908 2820 7936
rect 2700 6338 2728 7908
rect 2778 7848 2834 7857
rect 2778 7783 2834 7792
rect 2792 7546 2820 7783
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2884 7342 2912 10775
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2962 10024 3018 10033
rect 2962 9959 2964 9968
rect 3016 9959 3018 9968
rect 2964 9930 3016 9936
rect 3344 9738 3372 12406
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3436 10810 3464 12310
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3528 10742 3556 13903
rect 3608 13874 3660 13880
rect 3620 13569 3648 13874
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3620 12617 3648 12786
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3620 11558 3648 12378
rect 3712 11898 3740 19230
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3804 18358 3832 19110
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 3896 17746 3924 20216
rect 3884 17740 3936 17746
rect 3884 17682 3936 17688
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 3804 15366 3832 16186
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 12918 3832 13670
rect 3896 13462 3924 17478
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3804 11642 3832 12242
rect 3896 11762 3924 13262
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3712 11614 3832 11642
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3606 11384 3662 11393
rect 3712 11354 3740 11614
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3606 11319 3662 11328
rect 3700 11348 3752 11354
rect 3620 11286 3648 11319
rect 3700 11290 3752 11296
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3698 11248 3754 11257
rect 3698 11183 3754 11192
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3422 10568 3478 10577
rect 3422 10503 3478 10512
rect 3252 9710 3372 9738
rect 3252 9466 3280 9710
rect 3332 9648 3384 9654
rect 3330 9616 3332 9625
rect 3384 9616 3386 9625
rect 3436 9586 3464 10503
rect 3620 10266 3648 10950
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3606 10160 3662 10169
rect 3606 10095 3662 10104
rect 3514 9752 3570 9761
rect 3514 9687 3570 9696
rect 3330 9551 3386 9560
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3422 9480 3478 9489
rect 3252 9438 3372 9466
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3146 8936 3202 8945
rect 3146 8871 3202 8880
rect 3160 8362 3188 8871
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7449 3280 7686
rect 3238 7440 3294 7449
rect 3238 7375 3294 7384
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6458 2820 6734
rect 2884 6633 2912 6802
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 2870 6624 2926 6633
rect 2870 6559 2926 6568
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 3160 6361 3188 6695
rect 3252 6390 3280 6802
rect 3240 6384 3292 6390
rect 3146 6352 3202 6361
rect 2700 6310 2820 6338
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2792 4146 2820 6310
rect 3240 6326 3292 6332
rect 3146 6287 3202 6296
rect 2870 6216 2926 6225
rect 2870 6151 2926 6160
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 1214 4040 1270 4049
rect 388 4004 440 4010
rect 1214 3975 1270 3984
rect 388 3946 440 3952
rect 1228 3126 1256 3975
rect 2792 3738 2820 4082
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2884 3670 2912 6151
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3344 4826 3372 9438
rect 3422 9415 3424 9424
rect 3476 9415 3478 9424
rect 3424 9386 3476 9392
rect 3436 8498 3464 9386
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3528 5778 3556 9687
rect 3620 6458 3648 10095
rect 3712 6798 3740 11183
rect 3790 10840 3846 10849
rect 3790 10775 3792 10784
rect 3844 10775 3846 10784
rect 3792 10746 3844 10752
rect 3896 9738 3924 11494
rect 3988 11354 4016 20878
rect 4080 17678 4108 20998
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4172 20058 4200 20810
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4158 19000 4214 19009
rect 4158 18935 4214 18944
rect 4172 18834 4200 18935
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4068 17672 4120 17678
rect 4066 17640 4068 17649
rect 4120 17640 4122 17649
rect 4066 17575 4122 17584
rect 4264 17270 4292 23582
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4158 16008 4214 16017
rect 4158 15943 4214 15952
rect 4172 15162 4200 15943
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 14618 4200 14894
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4160 14340 4212 14346
rect 4160 14282 4212 14288
rect 4172 13938 4200 14282
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4066 12880 4122 12889
rect 4066 12815 4068 12824
rect 4120 12815 4122 12824
rect 4068 12786 4120 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4066 12472 4122 12481
rect 4066 12407 4068 12416
rect 4120 12407 4122 12416
rect 4068 12378 4120 12384
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4080 10266 4108 12271
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3804 9710 3924 9738
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3528 4826 3556 5578
rect 3804 5302 3832 9710
rect 3974 9616 4030 9625
rect 3884 9580 3936 9586
rect 3974 9551 4030 9560
rect 3884 9522 3936 9528
rect 3896 9382 3924 9522
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3896 9217 3924 9318
rect 3882 9208 3938 9217
rect 3882 9143 3938 9152
rect 3882 9072 3938 9081
rect 3882 9007 3938 9016
rect 3896 8106 3924 9007
rect 3988 8974 4016 9551
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3896 8078 4016 8106
rect 3988 6780 4016 8078
rect 3896 6752 4016 6780
rect 3896 5642 3924 6752
rect 4080 6458 4108 9930
rect 4172 9024 4200 12718
rect 4264 9654 4292 15438
rect 4356 15366 4384 21830
rect 4448 16182 4476 24822
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4540 22094 4568 23598
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4632 22409 4660 22578
rect 4618 22400 4674 22409
rect 4618 22335 4674 22344
rect 4540 22066 4660 22094
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 19514 4568 19722
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4434 15600 4490 15609
rect 4434 15535 4490 15544
rect 4344 15360 4396 15366
rect 4342 15328 4344 15337
rect 4396 15328 4398 15337
rect 4342 15263 4398 15272
rect 4448 15178 4476 15535
rect 4356 15150 4476 15178
rect 4356 13326 4384 15150
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4448 13977 4476 14214
rect 4434 13968 4490 13977
rect 4434 13903 4490 13912
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4434 13288 4490 13297
rect 4434 13223 4490 13232
rect 4448 13190 4476 13223
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4342 12336 4398 12345
rect 4342 12271 4398 12280
rect 4356 12102 4384 12271
rect 4344 12096 4396 12102
rect 4448 12073 4476 13126
rect 4344 12038 4396 12044
rect 4434 12064 4490 12073
rect 4434 11999 4490 12008
rect 4540 10266 4568 19246
rect 4632 17746 4660 22066
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4724 16590 4752 24278
rect 5276 22710 5304 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26330 7434 27000
rect 8022 26330 8078 27000
rect 6932 26302 7434 26330
rect 5460 23662 5488 26200
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23186 5580 23462
rect 6104 23186 6132 26200
rect 6276 25560 6328 25566
rect 6276 25502 6328 25508
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5172 22704 5224 22710
rect 5172 22646 5224 22652
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5184 21457 5212 22646
rect 5264 22500 5316 22506
rect 5264 22442 5316 22448
rect 5170 21448 5226 21457
rect 5170 21383 5226 21392
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4908 19514 4936 19790
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 17610 4844 18566
rect 4908 18154 4936 19450
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4896 17060 4948 17066
rect 4896 17002 4948 17008
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4710 15872 4766 15881
rect 4710 15807 4766 15816
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4632 13394 4660 14758
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4618 12744 4674 12753
rect 4618 12679 4674 12688
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4526 9888 4582 9897
rect 4526 9823 4582 9832
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4252 9512 4304 9518
rect 4250 9480 4252 9489
rect 4304 9480 4306 9489
rect 4250 9415 4306 9424
rect 4172 8996 4476 9024
rect 4250 8936 4306 8945
rect 4250 8871 4252 8880
rect 4304 8871 4306 8880
rect 4344 8900 4396 8906
rect 4252 8842 4304 8848
rect 4344 8842 4396 8848
rect 4356 8566 4384 8842
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4342 7712 4398 7721
rect 4342 7647 4398 7656
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6361 4200 6802
rect 4250 6488 4306 6497
rect 4250 6423 4306 6432
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 4158 6352 4214 6361
rect 4158 6287 4160 6296
rect 3988 5778 4016 6287
rect 4212 6287 4214 6296
rect 4160 6258 4212 6264
rect 4160 6112 4212 6118
rect 4158 6080 4160 6089
rect 4212 6080 4214 6089
rect 4158 6015 4214 6024
rect 4158 5808 4214 5817
rect 3976 5772 4028 5778
rect 4158 5743 4214 5752
rect 3976 5714 4028 5720
rect 4172 5710 4200 5743
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3804 4826 3832 5238
rect 4080 4826 4108 5306
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3330 4720 3386 4729
rect 3330 4655 3386 4664
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2872 3664 2924 3670
rect 1306 3632 1362 3641
rect 3344 3618 3372 4655
rect 4264 4622 4292 6423
rect 4356 6322 4384 7647
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4448 6186 4476 8996
rect 4540 7546 4568 9823
rect 4632 8566 4660 12679
rect 4724 11898 4752 15807
rect 4816 14482 4844 15982
rect 4908 15570 4936 17002
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4908 14482 4936 15506
rect 5000 15162 5028 21286
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18902 5120 19246
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5184 17921 5212 21383
rect 5276 20602 5304 22442
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5552 22166 5580 22374
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5644 21962 5672 22986
rect 5998 21992 6054 22001
rect 5632 21956 5684 21962
rect 5998 21927 6054 21936
rect 5632 21898 5684 21904
rect 5644 21865 5672 21898
rect 5908 21888 5960 21894
rect 5630 21856 5686 21865
rect 5908 21830 5960 21836
rect 5630 21791 5686 21800
rect 5448 21344 5500 21350
rect 5920 21321 5948 21830
rect 5448 21286 5500 21292
rect 5906 21312 5962 21321
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 18426 5304 18634
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5368 18193 5396 18770
rect 5460 18601 5488 21286
rect 5906 21247 5962 21256
rect 5814 21176 5870 21185
rect 5814 21111 5816 21120
rect 5868 21111 5870 21120
rect 5908 21140 5960 21146
rect 5816 21082 5868 21088
rect 5908 21082 5960 21088
rect 5920 20806 5948 21082
rect 6012 21078 6040 21927
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5920 20641 5948 20742
rect 5906 20632 5962 20641
rect 5906 20567 5962 20576
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5644 20346 5672 20402
rect 5908 20392 5960 20398
rect 5552 19258 5580 20334
rect 5644 20318 5856 20346
rect 5908 20334 5960 20340
rect 5828 20262 5856 20318
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5632 19780 5684 19786
rect 5632 19722 5684 19728
rect 5644 19378 5672 19722
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5552 19230 5672 19258
rect 5446 18592 5502 18601
rect 5446 18527 5502 18536
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5354 18184 5410 18193
rect 5354 18119 5410 18128
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5170 17912 5226 17921
rect 5170 17847 5226 17856
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4816 14362 4844 14418
rect 4816 14334 5028 14362
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4710 10160 4766 10169
rect 4710 10095 4766 10104
rect 4724 9178 4752 10095
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4816 8650 4844 14214
rect 5000 13870 5028 14334
rect 5092 14226 5120 16730
rect 5170 15736 5226 15745
rect 5170 15671 5226 15680
rect 5184 14414 5212 15671
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5092 14198 5212 14226
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 5092 13870 5120 13942
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4894 13696 4950 13705
rect 4894 13631 4950 13640
rect 4908 12442 4936 13631
rect 5092 13546 5120 13806
rect 5000 13518 5120 13546
rect 5000 13161 5028 13518
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4986 13152 5042 13161
rect 4986 13087 5042 13096
rect 5000 12918 5028 13087
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 5000 12322 5028 12854
rect 4908 12294 5028 12322
rect 4908 12073 4936 12294
rect 4988 12096 5040 12102
rect 4894 12064 4950 12073
rect 4988 12038 5040 12044
rect 4894 11999 4950 12008
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4908 9178 4936 11086
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4816 8634 4936 8650
rect 4804 8628 4936 8634
rect 4856 8622 4936 8628
rect 4804 8570 4856 8576
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4802 8528 4858 8537
rect 4802 8463 4858 8472
rect 4710 7984 4766 7993
rect 4710 7919 4766 7928
rect 4618 7576 4674 7585
rect 4528 7540 4580 7546
rect 4724 7546 4752 7919
rect 4618 7511 4674 7520
rect 4712 7540 4764 7546
rect 4528 7482 4580 7488
rect 4526 7304 4582 7313
rect 4526 7239 4582 7248
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4448 5114 4476 5238
rect 4540 5234 4568 7239
rect 4632 6458 4660 7511
rect 4712 7482 4764 7488
rect 4724 7342 4752 7482
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4816 7018 4844 8463
rect 4908 8378 4936 8622
rect 5000 8498 5028 12038
rect 5092 10538 5120 13398
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4908 8350 5028 8378
rect 4894 8256 4950 8265
rect 4894 8191 4950 8200
rect 4908 7886 4936 8191
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4724 6990 4844 7018
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5234 4660 5646
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4724 5114 4752 6990
rect 4448 5086 4752 5114
rect 4724 4690 4752 5086
rect 5000 5030 5028 8350
rect 5092 6730 5120 9590
rect 5184 9586 5212 14198
rect 5276 13705 5304 18022
rect 5552 17338 5580 18362
rect 5644 18086 5672 19230
rect 5736 18426 5764 20198
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5828 19446 5856 19654
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5644 17105 5672 17138
rect 5630 17096 5686 17105
rect 5630 17031 5686 17040
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5446 16552 5502 16561
rect 5446 16487 5502 16496
rect 5460 16454 5488 16487
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5552 15502 5580 16934
rect 5630 16280 5686 16289
rect 5630 16215 5632 16224
rect 5684 16215 5686 16224
rect 5632 16186 5684 16192
rect 5828 15881 5856 19246
rect 5920 18873 5948 20334
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6104 19666 6132 21422
rect 6196 20534 6224 21830
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 5906 18864 5962 18873
rect 5906 18799 5962 18808
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 5814 15872 5870 15881
rect 5814 15807 5870 15816
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5262 13696 5318 13705
rect 5262 13631 5318 13640
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5276 11762 5304 13398
rect 5368 12986 5396 14350
rect 5460 13326 5488 15302
rect 5644 14958 5672 15642
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5552 13938 5580 14282
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5644 13870 5672 14894
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14074 5856 14758
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5632 13864 5684 13870
rect 5538 13832 5594 13841
rect 5632 13806 5684 13812
rect 5538 13767 5594 13776
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5552 13138 5580 13767
rect 5828 13326 5856 14010
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5460 13110 5580 13138
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5368 12889 5396 12922
rect 5354 12880 5410 12889
rect 5354 12815 5410 12824
rect 5460 12306 5488 13110
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5552 12306 5580 12922
rect 5630 12336 5686 12345
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5540 12300 5592 12306
rect 5630 12271 5686 12280
rect 5540 12242 5592 12248
rect 5354 12064 5410 12073
rect 5354 11999 5410 12008
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5276 10810 5304 11018
rect 5368 11014 5396 11999
rect 5540 11688 5592 11694
rect 5460 11636 5540 11642
rect 5460 11630 5592 11636
rect 5460 11614 5580 11630
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5460 10606 5488 11614
rect 5538 10976 5594 10985
rect 5538 10911 5594 10920
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5552 10062 5580 10911
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5170 9072 5226 9081
rect 5170 9007 5226 9016
rect 5184 8974 5212 9007
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5184 8634 5212 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5276 7886 5304 9930
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5368 7546 5396 8910
rect 5460 8430 5488 9522
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5644 7834 5672 12271
rect 5736 11898 5764 13126
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5828 9908 5856 13126
rect 5920 10810 5948 18634
rect 6012 18222 6040 19654
rect 6104 19638 6224 19666
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6012 17921 6040 18022
rect 5998 17912 6054 17921
rect 5998 17847 6054 17856
rect 6012 15609 6040 17847
rect 6104 16794 6132 19450
rect 6196 18034 6224 19638
rect 6288 19553 6316 25502
rect 6644 25084 6696 25090
rect 6644 25026 6696 25032
rect 6458 24984 6514 24993
rect 6458 24919 6514 24928
rect 6472 22982 6500 24919
rect 6656 23526 6684 25026
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6460 22976 6512 22982
rect 6460 22918 6512 22924
rect 6458 22536 6514 22545
rect 6458 22471 6514 22480
rect 6472 22438 6500 22471
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6564 22386 6592 23462
rect 6748 22522 6776 26200
rect 6932 24290 6960 26302
rect 7378 26200 7434 26302
rect 7852 26302 8078 26330
rect 7378 25528 7434 25537
rect 7378 25463 7434 25472
rect 7104 24880 7156 24886
rect 7104 24822 7156 24828
rect 6840 24274 6960 24290
rect 6828 24268 6960 24274
rect 6880 24262 6960 24268
rect 6828 24210 6880 24216
rect 6828 23248 6880 23254
rect 6826 23216 6828 23225
rect 6880 23216 6882 23225
rect 6826 23151 6882 23160
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6918 22672 6974 22681
rect 6918 22607 6920 22616
rect 6972 22607 6974 22616
rect 6920 22578 6972 22584
rect 6748 22494 6960 22522
rect 6564 22358 6868 22386
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6552 20868 6604 20874
rect 6552 20810 6604 20816
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6274 19544 6330 19553
rect 6274 19479 6276 19488
rect 6328 19479 6330 19488
rect 6276 19450 6328 19456
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6288 19174 6316 19314
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6196 18006 6316 18034
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6196 16998 6224 17818
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6090 16280 6146 16289
rect 6090 16215 6146 16224
rect 5998 15600 6054 15609
rect 5998 15535 6054 15544
rect 5998 15056 6054 15065
rect 5998 14991 6000 15000
rect 6052 14991 6054 15000
rect 6000 14962 6052 14968
rect 6012 13530 6040 14962
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6012 12782 6040 13330
rect 6104 12918 6132 16215
rect 6196 15026 6224 16934
rect 6288 16674 6316 18006
rect 6380 17066 6408 20402
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 6366 16824 6422 16833
rect 6366 16759 6422 16768
rect 6380 16674 6408 16759
rect 6288 16646 6408 16674
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6196 13394 6224 13806
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6092 12912 6144 12918
rect 6090 12880 6092 12889
rect 6144 12880 6146 12889
rect 6196 12850 6224 13330
rect 6288 13258 6316 16458
rect 6380 16046 6408 16646
rect 6472 16454 6500 20538
rect 6564 19417 6592 20810
rect 6656 20398 6684 22170
rect 6840 22094 6868 22358
rect 6932 22166 6960 22494
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6748 22066 6868 22094
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6748 19938 6776 22066
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6932 21350 6960 21626
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 7024 21026 7052 23054
rect 7116 22710 7144 24822
rect 7392 24206 7420 25463
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7104 22704 7156 22710
rect 7104 22646 7156 22652
rect 7392 22574 7420 23054
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7392 22409 7420 22510
rect 7378 22400 7434 22409
rect 7378 22335 7434 22344
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 6932 20998 7052 21026
rect 6932 20482 6960 20998
rect 6932 20454 7052 20482
rect 6918 20360 6974 20369
rect 6918 20295 6974 20304
rect 6932 20058 6960 20295
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6748 19910 6960 19938
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6550 19408 6606 19417
rect 6656 19378 6684 19450
rect 6550 19343 6606 19352
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6748 17814 6776 19654
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6840 18834 6868 19314
rect 6932 19174 6960 19910
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6932 18766 6960 19110
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 18358 6960 18702
rect 7024 18465 7052 20454
rect 7010 18456 7066 18465
rect 7010 18391 7066 18400
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 17542 6592 17682
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6564 16250 6592 17478
rect 6656 17202 6684 17546
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6366 15600 6422 15609
rect 6564 15570 6592 15846
rect 6366 15535 6368 15544
rect 6420 15535 6422 15544
rect 6552 15564 6604 15570
rect 6368 15506 6420 15512
rect 6552 15506 6604 15512
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 13954 6408 14962
rect 6472 14074 6500 15370
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6380 13926 6500 13954
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6288 12889 6316 13194
rect 6274 12880 6330 12889
rect 6090 12815 6146 12824
rect 6184 12844 6236 12850
rect 6274 12815 6330 12824
rect 6184 12786 6236 12792
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12434 6040 12718
rect 6012 12406 6132 12434
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11898 6040 12038
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6104 11694 6132 12406
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6196 11336 6224 12786
rect 6380 12345 6408 13806
rect 6366 12336 6422 12345
rect 6366 12271 6368 12280
rect 6420 12271 6422 12280
rect 6368 12242 6420 12248
rect 6472 12186 6500 13926
rect 6564 12646 6592 15098
rect 6656 14006 6684 15846
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6012 11308 6224 11336
rect 6288 12158 6500 12186
rect 6552 12164 6604 12170
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10130 6040 11308
rect 6288 11234 6316 12158
rect 6552 12106 6604 12112
rect 6564 12073 6592 12106
rect 6550 12064 6606 12073
rect 6550 11999 6606 12008
rect 6656 11880 6684 13806
rect 6748 12850 6776 15574
rect 6840 13870 6868 17546
rect 6932 15026 6960 18022
rect 7012 17672 7064 17678
rect 7010 17640 7012 17649
rect 7064 17640 7066 17649
rect 7116 17626 7144 21354
rect 7208 18714 7236 21422
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7300 19378 7328 20266
rect 7484 19922 7512 24074
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7576 22098 7604 23598
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7576 21418 7604 22034
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7576 20398 7604 20810
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7392 19825 7420 19858
rect 7378 19816 7434 19825
rect 7378 19751 7434 19760
rect 7576 19446 7604 20334
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7208 18686 7328 18714
rect 7300 18630 7328 18686
rect 7288 18624 7340 18630
rect 7286 18592 7288 18601
rect 7340 18592 7342 18601
rect 7286 18527 7342 18536
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7116 17598 7236 17626
rect 7010 17575 7066 17584
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 16658 7144 17478
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7116 16153 7144 16458
rect 7102 16144 7158 16153
rect 7012 16108 7064 16114
rect 7102 16079 7158 16088
rect 7012 16050 7064 16056
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12918 6868 13262
rect 6932 12986 6960 13670
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 7024 12764 7052 16050
rect 7208 15994 7236 17598
rect 7300 17066 7328 18158
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7300 16658 7328 17002
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7392 16538 7420 18770
rect 7116 15966 7236 15994
rect 7300 16510 7420 16538
rect 7116 12832 7144 15966
rect 7300 14770 7328 16510
rect 7484 15366 7512 19382
rect 7576 19174 7604 19382
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7668 16454 7696 23666
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26330 10654 27000
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8128 23633 8156 23666
rect 8114 23624 8170 23633
rect 8114 23559 8170 23568
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 7840 22092 7892 22098
rect 7840 22034 7892 22040
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7656 16448 7708 16454
rect 7760 16425 7788 21898
rect 7852 21570 7880 22034
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8116 21616 8168 21622
rect 7852 21542 8064 21570
rect 8116 21558 8168 21564
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 7930 21448 7986 21457
rect 7852 21010 7880 21422
rect 7930 21383 7986 21392
rect 7944 21010 7972 21383
rect 8036 21146 8064 21542
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8128 21049 8156 21558
rect 8114 21040 8170 21049
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7932 21004 7984 21010
rect 8114 20975 8170 20984
rect 7932 20946 7984 20952
rect 7852 20330 7880 20946
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7840 20324 7892 20330
rect 7840 20266 7892 20272
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8220 20058 8248 20198
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 18834 7880 19926
rect 8312 19786 8340 21830
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 19961 8432 20742
rect 8390 19952 8446 19961
rect 8390 19887 8446 19896
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8312 19417 8340 19722
rect 8298 19408 8354 19417
rect 8298 19343 8354 19352
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 8300 18760 8352 18766
rect 8298 18728 8300 18737
rect 8352 18728 8354 18737
rect 8298 18663 8354 18672
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 18057 7880 18566
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8116 18352 8168 18358
rect 8036 18312 8116 18340
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7838 18048 7894 18057
rect 7838 17983 7894 17992
rect 7944 17921 7972 18090
rect 7930 17912 7986 17921
rect 7930 17847 7986 17856
rect 8036 17592 8064 18312
rect 8116 18294 8168 18300
rect 8206 18320 8262 18329
rect 8206 18255 8262 18264
rect 8114 18184 8170 18193
rect 8114 18119 8170 18128
rect 8128 17746 8156 18119
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7852 17564 8064 17592
rect 7852 16590 7880 17564
rect 8220 17542 8248 18255
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8404 17202 8432 18634
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8036 17054 8340 17082
rect 7932 16992 7984 16998
rect 7930 16960 7932 16969
rect 7984 16960 7986 16969
rect 7930 16895 7986 16904
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 8036 16436 8064 17054
rect 8312 16998 8340 17054
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8114 16688 8170 16697
rect 8114 16623 8116 16632
rect 8168 16623 8170 16632
rect 8116 16594 8168 16600
rect 7656 16390 7708 16396
rect 7746 16416 7802 16425
rect 7576 15706 7604 16390
rect 7746 16351 7802 16360
rect 7852 16408 8064 16436
rect 8220 16436 8248 16934
rect 8220 16408 8340 16436
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7562 15600 7618 15609
rect 7562 15535 7618 15544
rect 7472 15360 7524 15366
rect 7208 14742 7328 14770
rect 7392 15320 7472 15348
rect 7208 13530 7236 14742
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14074 7328 14214
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7208 13161 7236 13194
rect 7194 13152 7250 13161
rect 7194 13087 7250 13096
rect 7116 12804 7236 12832
rect 6932 12736 7052 12764
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6472 11852 6684 11880
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6104 11206 6316 11234
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5736 9880 5856 9908
rect 5736 7954 5764 9880
rect 5814 9752 5870 9761
rect 5814 9687 5870 9696
rect 5998 9752 6054 9761
rect 5998 9687 6054 9696
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5368 6390 5396 6734
rect 5552 6662 5580 7822
rect 5644 7806 5764 7834
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7342 5672 7686
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 6934 5672 7278
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5736 5370 5764 7806
rect 5828 7546 5856 9687
rect 6012 9654 6040 9687
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5906 9072 5962 9081
rect 5906 9007 5962 9016
rect 5920 8634 5948 9007
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 6012 6798 6040 8502
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 6458 6040 6734
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6104 5098 6132 11206
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10674 6316 10950
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6288 10470 6316 10610
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6274 9752 6330 9761
rect 6274 9687 6330 9696
rect 6288 9178 6316 9687
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6196 8634 6224 9114
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6288 8294 6316 8502
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7274 6224 7822
rect 6288 7546 6316 8230
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6288 7177 6316 7346
rect 6274 7168 6330 7177
rect 6274 7103 6330 7112
rect 6380 5846 6408 11630
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6472 5574 6500 11852
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6564 10266 6592 11698
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 10810 6684 11494
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6656 8480 6684 10406
rect 6748 8974 6776 12650
rect 6932 11354 6960 12736
rect 7208 12434 7236 12804
rect 7392 12434 7420 15320
rect 7472 15302 7524 15308
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 13530 7512 14758
rect 7576 14482 7604 15535
rect 7668 14550 7696 15982
rect 7760 15042 7788 15982
rect 7852 15502 7880 16408
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15706 7972 15914
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7944 15348 7972 15438
rect 7852 15320 7972 15348
rect 7852 15162 7880 15320
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7760 15014 7880 15042
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7576 13870 7604 14418
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 13394 7604 13806
rect 7564 13388 7616 13394
rect 7116 12406 7236 12434
rect 7300 12406 7420 12434
rect 7484 13348 7564 13376
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10010 7052 10950
rect 6840 9982 7052 10010
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6564 8452 6684 8480
rect 6736 8492 6788 8498
rect 6564 5778 6592 8452
rect 6736 8434 6788 8440
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6656 6798 6684 8298
rect 6748 8265 6776 8434
rect 6734 8256 6790 8265
rect 6734 8191 6790 8200
rect 6840 7834 6868 9982
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9466 6960 9862
rect 7012 9648 7064 9654
rect 7010 9616 7012 9625
rect 7064 9616 7066 9625
rect 7010 9551 7066 9560
rect 6932 9438 7052 9466
rect 6920 9376 6972 9382
rect 6918 9344 6920 9353
rect 6972 9344 6974 9353
rect 6918 9279 6974 9288
rect 7024 8090 7052 9438
rect 7116 9042 7144 12406
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7208 11626 7236 12310
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7300 11354 7328 12406
rect 7484 12186 7512 13348
rect 7564 13330 7616 13336
rect 7668 13274 7696 14486
rect 7760 14346 7788 14894
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7852 14226 7880 15014
rect 8220 14958 8248 15098
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 14385 8248 14418
rect 8206 14376 8262 14385
rect 8206 14311 8262 14320
rect 7760 14198 7880 14226
rect 7760 13938 7788 14198
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14074 8340 16408
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7576 13246 7696 13274
rect 7576 12306 7604 13246
rect 7760 12850 7788 13330
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12442 7696 12718
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7380 12164 7432 12170
rect 7484 12158 7604 12186
rect 7380 12106 7432 12112
rect 7392 12073 7420 12106
rect 7472 12096 7524 12102
rect 7378 12064 7434 12073
rect 7472 12038 7524 12044
rect 7378 11999 7434 12008
rect 7392 11830 7420 11999
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7392 11286 7420 11630
rect 7484 11558 7512 12038
rect 7576 11898 7604 12158
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7668 11778 7696 12106
rect 7576 11750 7696 11778
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7380 11280 7432 11286
rect 7286 11248 7342 11257
rect 7380 11222 7432 11228
rect 7286 11183 7342 11192
rect 7300 11150 7328 11183
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7208 7954 7236 10746
rect 7300 8650 7328 11086
rect 7392 10606 7420 11222
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7392 8838 7420 10367
rect 7484 10198 7512 11494
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7300 8622 7420 8650
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 6736 7812 6788 7818
rect 6840 7806 7236 7834
rect 6736 7754 6788 7760
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6254 6684 6734
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6748 5642 6776 7754
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7426 6960 7686
rect 6932 7398 7052 7426
rect 6828 7336 6880 7342
rect 6826 7304 6828 7313
rect 6920 7336 6972 7342
rect 6880 7304 6882 7313
rect 6920 7278 6972 7284
rect 6826 7239 6882 7248
rect 6932 7154 6960 7278
rect 7024 7206 7052 7398
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6840 7126 6960 7154
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6840 7002 6868 7126
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6840 6458 6868 6938
rect 6918 6896 6974 6905
rect 6918 6831 6974 6840
rect 6932 6662 6960 6831
rect 7116 6662 7144 7346
rect 7208 7188 7236 7806
rect 7392 7750 7420 8622
rect 7484 7818 7512 9046
rect 7576 8498 7604 11750
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7668 9178 7696 11630
rect 7760 10130 7788 12582
rect 7852 11150 7880 14010
rect 8404 13954 8432 16118
rect 8496 15978 8524 21626
rect 8588 20806 8616 22646
rect 8680 22574 8708 26200
rect 8852 26172 8904 26178
rect 8852 26114 8904 26120
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8864 21962 8892 26114
rect 9128 25016 9180 25022
rect 9128 24958 9180 24964
rect 8944 24132 8996 24138
rect 8944 24074 8996 24080
rect 8852 21956 8904 21962
rect 8852 21898 8904 21904
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8956 20482 8984 24074
rect 9140 23254 9168 24958
rect 9324 24342 9352 26200
rect 9864 25288 9916 25294
rect 9586 25256 9642 25265
rect 9864 25230 9916 25236
rect 9586 25191 9642 25200
rect 9772 25220 9824 25226
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9404 24336 9456 24342
rect 9404 24278 9456 24284
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9324 23497 9352 24142
rect 9416 23866 9444 24278
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9508 23526 9536 24006
rect 9496 23520 9548 23526
rect 9310 23488 9366 23497
rect 9496 23462 9548 23468
rect 9310 23423 9366 23432
rect 9128 23248 9180 23254
rect 9128 23190 9180 23196
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9310 22128 9366 22137
rect 9310 22063 9366 22072
rect 9324 21894 9352 22063
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9128 21616 9180 21622
rect 9128 21558 9180 21564
rect 9140 20534 9168 21558
rect 8772 20454 8984 20482
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8588 18193 8616 18770
rect 8574 18184 8630 18193
rect 8574 18119 8630 18128
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 8588 16114 8616 16458
rect 8680 16250 8708 16662
rect 8772 16590 8800 20454
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8864 19417 8892 20334
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8850 19408 8906 19417
rect 8850 19343 8906 19352
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16833 8892 17070
rect 8850 16824 8906 16833
rect 8850 16759 8906 16768
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8576 15904 8628 15910
rect 8482 15872 8538 15881
rect 8576 15846 8628 15852
rect 8482 15807 8538 15816
rect 8496 15570 8524 15807
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 15162 8524 15506
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8482 14648 8538 14657
rect 8482 14583 8484 14592
rect 8536 14583 8538 14592
rect 8484 14554 8536 14560
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8496 14278 8524 14418
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8588 14074 8616 15846
rect 8680 15570 8708 15982
rect 8772 15638 8800 16526
rect 8956 16402 8984 19450
rect 9140 19446 9168 20470
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 9232 19334 9260 21830
rect 9416 20262 9444 23054
rect 9494 22264 9550 22273
rect 9494 22199 9550 22208
rect 9508 20942 9536 22199
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9508 19990 9536 20334
rect 9496 19984 9548 19990
rect 9402 19952 9458 19961
rect 9496 19926 9548 19932
rect 9402 19887 9458 19896
rect 9416 19854 9444 19887
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9232 19306 9352 19334
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18970 9168 19110
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9048 18154 9076 18566
rect 9140 18290 9168 18906
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9140 17610 9168 18226
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 8864 16374 8984 16402
rect 8864 16250 8892 16374
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8312 13926 8432 13954
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 11286 7972 11766
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 8036 11218 8064 11834
rect 8114 11384 8170 11393
rect 8114 11319 8170 11328
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 8128 10996 8156 11319
rect 7852 10968 8156 10996
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7668 8430 7696 8910
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 8090 7604 8298
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7378 7440 7434 7449
rect 7378 7375 7380 7384
rect 7432 7375 7434 7384
rect 7472 7404 7524 7410
rect 7380 7346 7432 7352
rect 7472 7346 7524 7352
rect 7208 7160 7328 7188
rect 7300 7154 7328 7160
rect 7300 7126 7420 7154
rect 7194 7032 7250 7041
rect 7392 7002 7420 7126
rect 7194 6967 7196 6976
rect 7248 6967 7250 6976
rect 7380 6996 7432 7002
rect 7196 6938 7248 6944
rect 7380 6938 7432 6944
rect 6920 6656 6972 6662
rect 7104 6656 7156 6662
rect 6920 6598 6972 6604
rect 7010 6624 7066 6633
rect 7104 6598 7156 6604
rect 7010 6559 7066 6568
rect 6918 6488 6974 6497
rect 6828 6452 6880 6458
rect 6918 6423 6974 6432
rect 6828 6394 6880 6400
rect 6932 6118 6960 6423
rect 7024 6186 7052 6559
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7116 6118 7144 6598
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3436 3670 3464 4558
rect 3698 4448 3754 4457
rect 3698 4383 3754 4392
rect 3712 4146 3740 4383
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 2872 3606 2924 3612
rect 1306 3567 1308 3576
rect 1360 3567 1362 3576
rect 3252 3590 3372 3618
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 1308 3538 1360 3544
rect 3252 3194 3280 3590
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 1216 3120 1268 3126
rect 1216 3062 1268 3068
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 1308 2916 1360 2922
rect 1308 2858 1360 2864
rect 1320 2825 1348 2858
rect 1400 2848 1452 2854
rect 1306 2816 1362 2825
rect 1400 2790 1452 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1306 2751 1362 2760
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1216 2440 1268 2446
rect 1320 2417 1348 2450
rect 1216 2382 1268 2388
rect 1306 2408 1362 2417
rect 1228 2009 1256 2382
rect 1306 2343 1362 2352
rect 1308 2100 1360 2106
rect 1308 2042 1360 2048
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2042
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 1412 800 1440 2790
rect 2792 2446 2820 2790
rect 2884 2514 2912 2994
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3344 2310 3372 3470
rect 4080 3233 4108 3470
rect 4066 3224 4122 3233
rect 4066 3159 4122 3168
rect 7392 2990 7420 6938
rect 7484 3466 7512 7346
rect 7576 3738 7604 8026
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7668 6866 7696 7958
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7760 5846 7788 9862
rect 7852 9042 7880 10968
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10742 8340 13926
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8496 13326 8524 13738
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8680 13172 8708 15370
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 15094 8800 15302
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8772 14006 8800 15030
rect 8864 14385 8892 16050
rect 8956 14822 8984 16186
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8850 14376 8906 14385
rect 8850 14311 8906 14320
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8496 13144 8708 13172
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12102 8432 12582
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8404 10470 8432 11630
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 9994 8432 10406
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8404 9518 8432 9930
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8312 8537 8340 9454
rect 8298 8528 8354 8537
rect 8298 8463 8354 8472
rect 7840 8424 7892 8430
rect 8116 8424 8168 8430
rect 7840 8366 7892 8372
rect 8114 8392 8116 8401
rect 8168 8392 8170 8401
rect 7852 8294 7880 8366
rect 8114 8327 8170 8336
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 7410 7880 8230
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 7002 7880 7142
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5681 7880 6734
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7838 5672 7894 5681
rect 7838 5607 7894 5616
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 8312 4729 8340 8298
rect 8298 4720 8354 4729
rect 8298 4655 8354 4664
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2650 4384 2790
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 2106 3372 2246
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 4080 800 4108 2450
rect 6748 800 6776 2450
rect 8036 2310 8064 2926
rect 8312 2446 8340 3130
rect 8404 3058 8432 9454
rect 8496 8906 8524 13144
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8680 11354 8708 11562
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8772 10742 8800 11222
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8482 8256 8538 8265
rect 8482 8191 8538 8200
rect 8496 6730 8524 8191
rect 8588 8090 8616 10542
rect 8772 9654 8800 10678
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8680 8498 8708 8910
rect 8772 8498 8800 9046
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8680 7750 8708 8434
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8666 7576 8722 7585
rect 8666 7511 8722 7520
rect 8680 7410 8708 7511
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8496 6497 8524 6666
rect 8482 6488 8538 6497
rect 8680 6458 8708 7346
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8482 6423 8538 6432
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8772 3126 8800 7278
rect 8864 4554 8892 14214
rect 8956 14074 8984 14758
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8956 11762 8984 12174
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9048 10606 9076 17070
rect 9140 12238 9168 17546
rect 9232 17338 9260 18566
rect 9220 17332 9272 17338
rect 9324 17320 9352 19306
rect 9600 18873 9628 25191
rect 9772 25162 9824 25168
rect 9784 23610 9812 25162
rect 9876 23730 9904 25230
rect 9968 23798 9996 26200
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 9956 23792 10008 23798
rect 10060 23769 10088 24142
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 9956 23734 10008 23740
rect 10046 23760 10102 23769
rect 9864 23724 9916 23730
rect 10046 23695 10102 23704
rect 9864 23666 9916 23672
rect 9784 23582 9904 23610
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9692 22778 9720 22986
rect 9770 22944 9826 22953
rect 9770 22879 9826 22888
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9784 22642 9812 22879
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9876 22522 9904 23582
rect 9692 22494 9904 22522
rect 9692 20874 9720 22494
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9784 22098 9812 22170
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9956 22094 10008 22098
rect 10152 22094 10180 23802
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 9956 22092 10180 22094
rect 10008 22066 10180 22092
rect 9956 22034 10008 22040
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9784 19514 9812 21490
rect 9968 20641 9996 22034
rect 9954 20632 10010 20641
rect 9954 20567 10010 20576
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9586 18864 9642 18873
rect 9586 18799 9642 18808
rect 9678 18728 9734 18737
rect 9404 18692 9456 18698
rect 9678 18663 9734 18672
rect 9772 18692 9824 18698
rect 9404 18634 9456 18640
rect 9416 18290 9444 18634
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9404 17332 9456 17338
rect 9324 17292 9404 17320
rect 9220 17274 9272 17280
rect 9404 17274 9456 17280
rect 9416 16833 9444 17274
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 15586 9260 16390
rect 9416 16250 9444 16662
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9416 16017 9444 16050
rect 9402 16008 9458 16017
rect 9402 15943 9458 15952
rect 9508 15910 9536 18566
rect 9692 18358 9720 18663
rect 9772 18634 9824 18640
rect 9784 18601 9812 18634
rect 9770 18592 9826 18601
rect 9770 18527 9826 18536
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9588 18148 9640 18154
rect 9640 18108 9720 18136
rect 9588 18090 9640 18096
rect 9586 18048 9642 18057
rect 9692 18034 9720 18108
rect 9692 18006 9812 18034
rect 9586 17983 9642 17992
rect 9496 15904 9548 15910
rect 9600 15881 9628 17983
rect 9678 17912 9734 17921
rect 9784 17898 9812 18006
rect 9734 17870 9812 17898
rect 9678 17847 9734 17856
rect 9876 17610 9904 20198
rect 9968 19922 9996 20266
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17338 9720 17478
rect 9968 17354 9996 19450
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9876 17326 9996 17354
rect 9692 16794 9720 17274
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9784 16658 9812 16934
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9496 15846 9548 15852
rect 9586 15872 9642 15881
rect 9586 15807 9642 15816
rect 9416 15706 9674 15722
rect 9404 15700 9686 15706
rect 9456 15694 9634 15700
rect 9404 15642 9456 15648
rect 9634 15642 9686 15648
rect 9784 15638 9812 16594
rect 9876 16522 9904 17326
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9968 16425 9996 17138
rect 9954 16416 10010 16425
rect 9954 16351 10010 16360
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9772 15632 9824 15638
rect 9232 15570 9674 15586
rect 9772 15574 9824 15580
rect 9232 15564 9686 15570
rect 9232 15558 9634 15564
rect 9634 15506 9686 15512
rect 9876 15502 9904 15846
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9404 15428 9456 15434
rect 9588 15428 9640 15434
rect 9456 15388 9588 15416
rect 9404 15370 9456 15376
rect 9588 15370 9640 15376
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9496 15088 9548 15094
rect 9232 15048 9496 15076
rect 9232 14550 9260 15048
rect 9496 15030 9548 15036
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9600 14278 9628 14758
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11830 9168 12174
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8956 9654 8984 9687
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8956 8974 8984 9590
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8956 4010 8984 7346
rect 9048 5914 9076 8774
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9140 5710 9168 10474
rect 9232 7886 9260 13126
rect 9324 12986 9352 13806
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9324 12306 9352 12922
rect 9416 12434 9444 13126
rect 9508 12850 9536 13942
rect 9588 13864 9640 13870
rect 9586 13832 9588 13841
rect 9640 13832 9642 13841
rect 9586 13767 9642 13776
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9416 12406 9536 12434
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9324 9722 9352 11154
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9416 8566 9444 9930
rect 9404 8560 9456 8566
rect 9310 8528 9366 8537
rect 9404 8502 9456 8508
rect 9310 8463 9366 8472
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9324 5914 9352 8463
rect 9402 7984 9458 7993
rect 9402 7919 9404 7928
rect 9456 7919 9458 7928
rect 9404 7890 9456 7896
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6322 9444 6734
rect 9508 6322 9536 12406
rect 9600 10674 9628 13670
rect 9692 11150 9720 15302
rect 9770 14648 9826 14657
rect 9770 14583 9826 14592
rect 9784 14550 9812 14583
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9876 14482 9904 15302
rect 9968 15094 9996 16351
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 11529 9812 13330
rect 9770 11520 9826 11529
rect 9770 11455 9826 11464
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9772 11008 9824 11014
rect 9770 10976 9772 10985
rect 9824 10976 9826 10985
rect 9692 10934 9770 10962
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9600 9110 9628 10610
rect 9692 9466 9720 10934
rect 9770 10911 9826 10920
rect 9876 10130 9904 14214
rect 9968 11286 9996 14758
rect 10060 13705 10088 19722
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10152 19281 10180 19314
rect 10138 19272 10194 19281
rect 10138 19207 10194 19216
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10152 16522 10180 18770
rect 10244 17377 10272 23598
rect 10704 22710 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 11060 25424 11112 25430
rect 11060 25366 11112 25372
rect 11072 22817 11100 25366
rect 11150 23896 11206 23905
rect 11150 23831 11206 23840
rect 11164 23254 11192 23831
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11058 22808 11114 22817
rect 11058 22743 11060 22752
rect 11112 22743 11114 22752
rect 11060 22714 11112 22720
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10692 22160 10744 22166
rect 10876 22160 10928 22166
rect 10744 22120 10876 22148
rect 10692 22102 10744 22108
rect 10876 22102 10928 22108
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10600 22024 10652 22030
rect 10876 22024 10928 22030
rect 10652 22001 10732 22012
rect 10652 21992 10746 22001
rect 10652 21984 10690 21992
rect 10600 21966 10652 21972
rect 10520 21729 10548 21966
rect 10876 21966 10928 21972
rect 10690 21927 10746 21936
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10506 21720 10562 21729
rect 10506 21655 10562 21664
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10336 18834 10364 21422
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10506 21312 10562 21321
rect 10428 21049 10456 21286
rect 10506 21247 10562 21256
rect 10414 21040 10470 21049
rect 10414 20975 10470 20984
rect 10520 20641 10548 21247
rect 10612 20777 10640 21830
rect 10888 21690 10916 21966
rect 10980 21690 11008 22510
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22273 11100 22374
rect 11058 22264 11114 22273
rect 11164 22234 11192 22510
rect 11058 22199 11114 22208
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11060 21956 11112 21962
rect 11060 21898 11112 21904
rect 11072 21729 11100 21898
rect 11058 21720 11114 21729
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10968 21684 11020 21690
rect 11058 21655 11114 21664
rect 10968 21626 11020 21632
rect 10876 21480 10928 21486
rect 10968 21480 11020 21486
rect 10876 21422 10928 21428
rect 10966 21448 10968 21457
rect 11020 21448 11022 21457
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10598 20768 10654 20777
rect 10598 20703 10654 20712
rect 10506 20632 10562 20641
rect 10506 20567 10562 20576
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10704 19689 10732 20402
rect 10796 20210 10824 21354
rect 10888 20398 10916 21422
rect 10966 21383 11022 21392
rect 11164 21321 11192 22170
rect 11256 22098 11284 26200
rect 11796 25764 11848 25770
rect 11796 25706 11848 25712
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 23050 11744 24006
rect 11428 23044 11480 23050
rect 11428 22986 11480 22992
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11348 22234 11376 22578
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11440 21350 11468 22986
rect 11808 22930 11836 25706
rect 11716 22902 11836 22930
rect 11716 21865 11744 22902
rect 11794 22808 11850 22817
rect 11794 22743 11850 22752
rect 11808 22710 11836 22743
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11702 21856 11758 21865
rect 11702 21791 11758 21800
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11428 21344 11480 21350
rect 11150 21312 11206 21321
rect 11428 21286 11480 21292
rect 11150 21247 11206 21256
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 11060 20256 11112 20262
rect 10796 20182 10916 20210
rect 11060 20198 11112 20204
rect 10690 19680 10746 19689
rect 10690 19615 10746 19624
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10428 18970 10456 19246
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18193 10364 18566
rect 10322 18184 10378 18193
rect 10322 18119 10378 18128
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10230 17368 10286 17377
rect 10336 17338 10364 17818
rect 10428 17762 10456 18702
rect 10520 17882 10548 19246
rect 10704 19145 10732 19615
rect 10888 19334 10916 20182
rect 11072 19786 11100 20198
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 11072 19446 11100 19722
rect 11060 19440 11112 19446
rect 11164 19417 11192 20742
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11060 19382 11112 19388
rect 11150 19408 11206 19417
rect 11150 19343 11206 19352
rect 10888 19306 11008 19334
rect 10784 19168 10836 19174
rect 10690 19136 10746 19145
rect 10784 19110 10836 19116
rect 10874 19136 10930 19145
rect 10690 19071 10746 19080
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10612 18737 10640 18838
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 10598 18728 10654 18737
rect 10598 18663 10654 18672
rect 10704 18329 10732 18770
rect 10796 18578 10824 19110
rect 10874 19071 10930 19080
rect 10888 18834 10916 19071
rect 10980 18902 11008 19306
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 11060 18624 11112 18630
rect 10796 18550 11008 18578
rect 11060 18566 11112 18572
rect 10690 18320 10746 18329
rect 10690 18255 10746 18264
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10612 18057 10640 18158
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10598 18048 10654 18057
rect 10598 17983 10654 17992
rect 10888 17921 10916 18090
rect 10874 17912 10930 17921
rect 10508 17876 10560 17882
rect 10874 17847 10930 17856
rect 10508 17818 10560 17824
rect 10428 17734 10548 17762
rect 10230 17303 10286 17312
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10336 17134 10364 17274
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10152 16114 10180 16458
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10152 15201 10180 16050
rect 10138 15192 10194 15201
rect 10138 15127 10194 15136
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10152 14482 10180 15030
rect 10244 14482 10272 17070
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10138 14376 10194 14385
rect 10138 14311 10194 14320
rect 10046 13696 10102 13705
rect 10046 13631 10102 13640
rect 10152 13274 10180 14311
rect 10336 14074 10364 15506
rect 10428 15502 10456 16934
rect 10520 16182 10548 17734
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10612 16833 10640 17478
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10598 16824 10654 16833
rect 10598 16759 10654 16768
rect 10600 16584 10652 16590
rect 10704 16572 10732 17002
rect 10652 16544 10732 16572
rect 10600 16526 10652 16532
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10520 16017 10548 16118
rect 10704 16046 10732 16544
rect 10600 16040 10652 16046
rect 10506 16008 10562 16017
rect 10600 15982 10652 15988
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10506 15943 10562 15952
rect 10612 15910 10640 15982
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10520 14822 10548 15642
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 14958 10640 15506
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10612 14498 10640 14894
rect 10704 14793 10732 14962
rect 10690 14784 10746 14793
rect 10690 14719 10746 14728
rect 10428 14470 10640 14498
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10244 13870 10272 14010
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10336 13734 10364 14010
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10060 13246 10180 13274
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9876 9761 9904 9930
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9876 9518 9904 9687
rect 9864 9512 9916 9518
rect 9692 9438 9812 9466
rect 9864 9454 9916 9460
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8566 9628 8842
rect 9692 8634 9720 9007
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9692 8090 9720 8570
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9678 7032 9734 7041
rect 9678 6967 9734 6976
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9692 6254 9720 6967
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9784 5914 9812 9438
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8634 9904 8842
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 8265 9904 8366
rect 9862 8256 9918 8265
rect 9862 8191 9918 8200
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9876 8022 9904 8055
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7449 9904 7822
rect 9862 7440 9918 7449
rect 9862 7375 9918 7384
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9968 4758 9996 11086
rect 10060 10538 10088 13246
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 8129 10088 9318
rect 10152 9178 10180 13126
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10244 12850 10272 12951
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10046 8120 10102 8129
rect 10046 8055 10102 8064
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9956 4752 10008 4758
rect 9956 4694 10008 4700
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8392 3052 8444 3058
rect 10060 3040 10088 7686
rect 10152 4826 10180 8910
rect 10244 7274 10272 12174
rect 10336 9926 10364 13126
rect 10428 12918 10456 14470
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10612 12986 10640 14350
rect 10796 13818 10824 17478
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16114 10916 16934
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10980 15881 11008 18550
rect 11072 17513 11100 18566
rect 11164 18329 11192 19110
rect 11256 18816 11284 20470
rect 11440 20262 11468 21286
rect 11532 21010 11560 21354
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11624 20210 11652 21490
rect 11716 20534 11744 21791
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11808 20890 11836 21558
rect 11900 21010 11928 26200
rect 12440 25968 12492 25974
rect 12440 25910 12492 25916
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12084 24449 12112 25298
rect 12070 24440 12126 24449
rect 12070 24375 12126 24384
rect 11978 24304 12034 24313
rect 11978 24239 12034 24248
rect 11992 23662 12020 24239
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12084 23050 12112 24375
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11808 20862 11928 20890
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11348 19718 11376 19926
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11440 19446 11468 20198
rect 11624 20182 11836 20210
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11518 19952 11574 19961
rect 11518 19887 11574 19896
rect 11532 19553 11560 19887
rect 11624 19854 11652 19994
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11518 19544 11574 19553
rect 11518 19479 11574 19488
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11440 19334 11468 19382
rect 11348 19306 11468 19334
rect 11348 18986 11376 19306
rect 11532 19258 11560 19479
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11440 19230 11560 19258
rect 11440 19174 11468 19230
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11348 18958 11560 18986
rect 11532 18816 11560 18958
rect 11612 18896 11664 18902
rect 11256 18788 11376 18816
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11150 18320 11206 18329
rect 11150 18255 11206 18264
rect 11150 18048 11206 18057
rect 11150 17983 11206 17992
rect 11058 17504 11114 17513
rect 11058 17439 11114 17448
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16289 11100 16390
rect 11058 16280 11114 16289
rect 11058 16215 11114 16224
rect 11060 15904 11112 15910
rect 10966 15872 11022 15881
rect 11060 15846 11112 15852
rect 10966 15807 11022 15816
rect 10966 14784 11022 14793
rect 10966 14719 11022 14728
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10704 13790 10824 13818
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11354 10456 12106
rect 10520 11898 10548 12854
rect 10704 12434 10732 13790
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10612 12406 10732 12434
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10506 11792 10562 11801
rect 10506 11727 10562 11736
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10520 11257 10548 11727
rect 10506 11248 10562 11257
rect 10506 11183 10562 11192
rect 10612 10826 10640 12406
rect 10796 12186 10824 13262
rect 10888 12918 10916 14350
rect 10980 13954 11008 14719
rect 11072 14278 11100 15846
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10980 13926 11100 13954
rect 10966 13832 11022 13841
rect 10966 13767 10968 13776
rect 11020 13767 11022 13776
rect 10968 13738 11020 13744
rect 11072 13462 11100 13926
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 11164 12764 11192 17983
rect 10888 12736 11192 12764
rect 10888 12442 10916 12736
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12442 11008 12582
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10704 12158 10824 12186
rect 10704 11626 10732 12158
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10520 10798 10640 10826
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10322 9616 10378 9625
rect 10322 9551 10378 9560
rect 10336 9042 10364 9551
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10322 8800 10378 8809
rect 10322 8735 10378 8744
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10336 6866 10364 8735
rect 10428 8634 10456 10406
rect 10520 9897 10548 10798
rect 10598 10704 10654 10713
rect 10598 10639 10654 10648
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8566 10548 9658
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10612 8378 10640 10639
rect 10690 9752 10746 9761
rect 10690 9687 10746 9696
rect 10704 9654 10732 9687
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 10690 9072 10746 9081
rect 10690 9007 10746 9016
rect 10704 8974 10732 9007
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10428 8350 10640 8378
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10428 6322 10456 8350
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10612 7562 10640 7890
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10520 7534 10640 7562
rect 10520 7410 10548 7534
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10506 6760 10562 6769
rect 10506 6695 10508 6704
rect 10560 6695 10562 6704
rect 10508 6666 10560 6672
rect 10612 6458 10640 7346
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10704 5574 10732 7822
rect 10796 7546 10824 12038
rect 10888 10742 10916 12242
rect 10980 10810 11008 12378
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10876 10736 10928 10742
rect 11072 10690 11100 11766
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 10849 11192 11154
rect 11150 10840 11206 10849
rect 11150 10775 11206 10784
rect 10876 10678 10928 10684
rect 10980 10662 11100 10690
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9722 10916 9862
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 8974 10916 9318
rect 10980 9081 11008 10662
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9722 11192 9862
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 10966 9072 11022 9081
rect 10966 9007 11022 9016
rect 10876 8968 10928 8974
rect 10928 8928 11008 8956
rect 10876 8910 10928 8916
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10888 6882 10916 8774
rect 10980 7562 11008 8928
rect 11058 8664 11114 8673
rect 11058 8599 11060 8608
rect 11112 8599 11114 8608
rect 11060 8570 11112 8576
rect 11164 8537 11192 9454
rect 11150 8528 11206 8537
rect 11150 8463 11206 8472
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7750 11100 8298
rect 11256 7886 11284 18566
rect 11348 17746 11376 18788
rect 11440 18788 11560 18816
rect 11610 18864 11612 18873
rect 11664 18864 11666 18873
rect 11610 18799 11666 18808
rect 11440 18086 11468 18788
rect 11610 18456 11666 18465
rect 11610 18391 11666 18400
rect 11518 18320 11574 18329
rect 11518 18255 11574 18264
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11348 13326 11376 17546
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11440 16522 11468 17138
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11426 16280 11482 16289
rect 11426 16215 11482 16224
rect 11440 15638 11468 16215
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11532 15484 11560 18255
rect 11624 18222 11652 18391
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11716 17746 11744 19314
rect 11808 19145 11836 20182
rect 11794 19136 11850 19145
rect 11794 19071 11850 19080
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11808 18465 11836 18634
rect 11794 18456 11850 18465
rect 11794 18391 11850 18400
rect 11796 18352 11848 18358
rect 11794 18320 11796 18329
rect 11848 18320 11850 18329
rect 11794 18255 11850 18264
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11624 15910 11652 17682
rect 11716 16114 11744 17682
rect 11796 16992 11848 16998
rect 11794 16960 11796 16969
rect 11848 16960 11850 16969
rect 11794 16895 11850 16904
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11808 16425 11836 16526
rect 11794 16416 11850 16425
rect 11794 16351 11850 16360
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11612 15496 11664 15502
rect 11532 15456 11612 15484
rect 11664 15456 11744 15484
rect 11612 15438 11664 15444
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11440 14113 11468 15370
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11426 14104 11482 14113
rect 11426 14039 11482 14048
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 8838 11376 12582
rect 11532 12434 11560 15302
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14074 11652 14962
rect 11716 14618 11744 15456
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11716 14521 11744 14554
rect 11702 14512 11758 14521
rect 11702 14447 11758 14456
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11624 13977 11652 14010
rect 11610 13968 11666 13977
rect 11610 13903 11666 13912
rect 11716 13462 11744 14214
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11440 12406 11560 12434
rect 11440 9353 11468 12406
rect 11716 11880 11744 13194
rect 11808 12617 11836 15846
rect 11900 12986 11928 20862
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11992 20505 12020 20538
rect 11978 20496 12034 20505
rect 11978 20431 12034 20440
rect 11978 19952 12034 19961
rect 11978 19887 12034 19896
rect 11992 19334 12020 19887
rect 11992 19310 12112 19334
rect 11992 19306 12124 19310
rect 12072 19304 12124 19306
rect 12176 19281 12204 21422
rect 12268 20806 12296 25638
rect 12452 23202 12480 25910
rect 12544 23798 12572 26200
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12360 23174 12480 23202
rect 12532 23180 12584 23186
rect 12360 22030 12388 23174
rect 12532 23122 12584 23128
rect 12544 22778 12572 23122
rect 12636 23089 12664 24142
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12636 22778 12664 22918
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12544 22094 12572 22714
rect 12728 22710 12756 22918
rect 13174 22808 13230 22817
rect 13174 22743 13230 22752
rect 12716 22704 12768 22710
rect 12716 22646 12768 22652
rect 12728 22094 12756 22646
rect 13188 22545 13216 22743
rect 13174 22536 13230 22545
rect 13174 22471 13230 22480
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22098 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15566 26208 15622 26217
rect 13634 26072 13690 26081
rect 13634 26007 13690 26016
rect 13544 25492 13596 25498
rect 13544 25434 13596 25440
rect 12452 22066 12572 22094
rect 12636 22066 12756 22094
rect 13360 22092 13412 22098
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12360 21593 12388 21966
rect 12452 21690 12480 22066
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12532 21616 12584 21622
rect 12346 21584 12402 21593
rect 12346 21519 12402 21528
rect 12530 21584 12532 21593
rect 12584 21584 12586 21593
rect 12530 21519 12586 21528
rect 12348 20936 12400 20942
rect 12346 20904 12348 20913
rect 12400 20904 12402 20913
rect 12346 20839 12402 20848
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12268 19904 12296 20742
rect 12360 20262 12388 20742
rect 12530 20496 12586 20505
rect 12530 20431 12586 20440
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12544 19961 12572 20431
rect 12530 19952 12586 19961
rect 12268 19876 12480 19904
rect 12530 19887 12586 19896
rect 12346 19816 12402 19825
rect 12346 19751 12348 19760
rect 12400 19751 12402 19760
rect 12348 19722 12400 19728
rect 12256 19712 12308 19718
rect 12452 19666 12480 19876
rect 12256 19654 12308 19660
rect 12072 19246 12124 19252
rect 12162 19272 12218 19281
rect 12162 19207 12218 19216
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18630 12020 18702
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18465 12112 18566
rect 12070 18456 12126 18465
rect 12070 18391 12126 18400
rect 12176 18136 12204 18770
rect 12268 18714 12296 19654
rect 12360 19638 12480 19666
rect 12360 19009 12388 19638
rect 12636 19530 12664 22066
rect 13360 22034 13412 22040
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21729 13124 21966
rect 13358 21856 13414 21865
rect 13358 21791 13414 21800
rect 13082 21720 13138 21729
rect 13082 21655 13138 21664
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12728 20942 12756 21354
rect 12820 21185 12848 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12806 21176 12862 21185
rect 12950 21179 13258 21188
rect 12806 21111 12862 21120
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12716 20256 12768 20262
rect 12820 20233 12848 20470
rect 13372 20398 13400 21791
rect 13556 21486 13584 25434
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13450 21176 13506 21185
rect 13450 21111 13506 21120
rect 13464 21010 13492 21111
rect 13556 21078 13584 21286
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13648 20534 13676 26007
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13740 24177 13768 24647
rect 13726 24168 13782 24177
rect 13832 24138 13860 26200
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14292 24342 14320 24754
rect 14476 24562 14504 26200
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 14830 24848 14886 24857
rect 14830 24783 14886 24792
rect 14384 24534 14504 24562
rect 14554 24576 14610 24585
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14384 24274 14412 24534
rect 14554 24511 14610 24520
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14464 24200 14516 24206
rect 14568 24177 14596 24511
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14464 24142 14516 24148
rect 14554 24168 14610 24177
rect 13726 24103 13782 24112
rect 13820 24132 13872 24138
rect 13740 23730 13768 24103
rect 13820 24074 13872 24080
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13832 22642 13860 22986
rect 13820 22636 13872 22642
rect 13872 22596 13952 22624
rect 13820 22578 13872 22584
rect 13924 22166 13952 22596
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 13912 22160 13964 22166
rect 13818 22128 13874 22137
rect 13912 22102 13964 22108
rect 13818 22063 13874 22072
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 13740 20466 13768 21558
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13360 20392 13412 20398
rect 13358 20360 13360 20369
rect 13412 20360 13414 20369
rect 13358 20295 13414 20304
rect 12716 20198 12768 20204
rect 12806 20224 12862 20233
rect 12452 19502 12664 19530
rect 12346 19000 12402 19009
rect 12452 18970 12480 19502
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12346 18935 12402 18944
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12268 18686 12388 18714
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 11992 18108 12204 18136
rect 11992 15910 12020 18108
rect 12268 17762 12296 18566
rect 12360 18057 12388 18686
rect 12544 18290 12572 18838
rect 12636 18766 12664 19246
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12440 18080 12492 18086
rect 12346 18048 12402 18057
rect 12440 18022 12492 18028
rect 12346 17983 12402 17992
rect 12176 17734 12296 17762
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12084 16794 12112 17138
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11978 15192 12034 15201
rect 11978 15127 12034 15136
rect 11992 14550 12020 15127
rect 11980 14544 12032 14550
rect 11978 14512 11980 14521
rect 12032 14512 12034 14521
rect 11978 14447 12034 14456
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13394 12020 14350
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11978 12880 12034 12889
rect 11978 12815 12034 12824
rect 11794 12608 11850 12617
rect 11794 12543 11850 12552
rect 11794 12200 11850 12209
rect 11794 12135 11850 12144
rect 11808 12102 11836 12135
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11898 11928 12038
rect 11992 11937 12020 12815
rect 12084 12374 12112 16526
rect 12176 15586 12204 17734
rect 12452 17610 12480 18022
rect 12440 17604 12492 17610
rect 12360 17564 12440 17592
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12268 16182 12296 16730
rect 12360 16289 12388 17564
rect 12440 17546 12492 17552
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 12452 17066 12480 17439
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12346 16280 12402 16289
rect 12346 16215 12402 16224
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12452 15745 12480 16458
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12544 15609 12572 17002
rect 12636 16658 12664 17070
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12530 15600 12586 15609
rect 12176 15558 12296 15586
rect 12162 15464 12218 15473
rect 12162 15399 12218 15408
rect 12176 15366 12204 15399
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12268 15144 12296 15558
rect 12530 15535 12586 15544
rect 12636 15450 12664 16390
rect 12544 15422 12664 15450
rect 12440 15156 12492 15162
rect 12268 15116 12440 15144
rect 12440 15098 12492 15104
rect 12254 14512 12310 14521
rect 12544 14498 12572 15422
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12254 14447 12310 14456
rect 12452 14470 12572 14498
rect 12162 13968 12218 13977
rect 12162 13903 12164 13912
rect 12216 13903 12218 13912
rect 12164 13874 12216 13880
rect 12268 13512 12296 14447
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12176 13484 12296 13512
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 11978 11928 12034 11937
rect 11532 11852 11744 11880
rect 11888 11892 11940 11898
rect 11426 9344 11482 9353
rect 11426 9279 11482 9288
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11334 8664 11390 8673
rect 11334 8599 11336 8608
rect 11388 8599 11390 8608
rect 11336 8570 11388 8576
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10980 7546 11100 7562
rect 10980 7540 11112 7546
rect 10980 7534 11060 7540
rect 11060 7482 11112 7488
rect 11348 7449 11376 7958
rect 11334 7440 11390 7449
rect 11334 7375 11390 7384
rect 10796 6854 10916 6882
rect 10796 6662 10824 6854
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10784 6656 10836 6662
rect 10888 6633 10916 6666
rect 10784 6598 10836 6604
rect 10874 6624 10930 6633
rect 10874 6559 10930 6568
rect 11440 6458 11468 8502
rect 11532 7342 11560 11852
rect 11978 11863 12034 11872
rect 11888 11834 11940 11840
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11716 11098 11744 11727
rect 11624 10674 11652 11086
rect 11716 11082 11836 11098
rect 11716 11076 11848 11082
rect 11716 11070 11796 11076
rect 11716 10810 11744 11070
rect 11796 11018 11848 11024
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 9994 11652 10610
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11624 9586 11652 9930
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11716 9042 11744 9386
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11808 8922 11836 9930
rect 11716 8894 11836 8922
rect 11610 8664 11666 8673
rect 11610 8599 11612 8608
rect 11664 8599 11666 8608
rect 11612 8570 11664 8576
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11624 6798 11652 8298
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11716 6322 11744 8894
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 6798 11836 8774
rect 11900 6866 11928 11018
rect 11992 10810 12020 11863
rect 12070 11520 12126 11529
rect 12070 11455 12126 11464
rect 12084 10810 12112 11455
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11992 10538 12020 10746
rect 12176 10690 12204 13484
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 11694 12296 13330
rect 12360 12714 12388 13738
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 12452 12458 12480 14470
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12360 12430 12480 12458
rect 12360 12102 12388 12430
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12256 11688 12308 11694
rect 12452 11642 12480 12038
rect 12256 11630 12308 11636
rect 12360 11614 12480 11642
rect 12256 11552 12308 11558
rect 12360 11506 12388 11614
rect 12308 11500 12388 11506
rect 12256 11494 12388 11500
rect 12268 11478 12388 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12084 10662 12204 10690
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 9654 12020 9862
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11992 6254 12020 9454
rect 12084 7546 12112 10662
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 9994 12204 10406
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12176 9897 12204 9930
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12268 9738 12296 11154
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12176 9710 12296 9738
rect 12176 8906 12204 9710
rect 12360 9518 12388 10746
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8786 12296 8842
rect 12176 8758 12296 8786
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12176 7206 12204 8758
rect 12360 8362 12388 9454
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12346 8120 12402 8129
rect 12346 8055 12348 8064
rect 12400 8055 12402 8064
rect 12348 8026 12400 8032
rect 12452 7818 12480 11290
rect 12544 8838 12572 14282
rect 12636 12102 12664 15302
rect 12728 14385 12756 20198
rect 12806 20159 12862 20168
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12990 19816 13046 19825
rect 12808 19780 12860 19786
rect 12990 19751 13046 19760
rect 12808 19722 12860 19728
rect 12820 19334 12848 19722
rect 13004 19718 13032 19751
rect 13556 19718 13584 20402
rect 13740 19990 13768 20402
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 12820 19306 13124 19334
rect 13096 19174 13124 19306
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18465 13400 19654
rect 13358 18456 13414 18465
rect 13358 18391 13414 18400
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12992 18216 13044 18222
rect 12990 18184 12992 18193
rect 13044 18184 13046 18193
rect 12808 18148 12860 18154
rect 13096 18170 13124 18226
rect 13096 18142 13400 18170
rect 13464 18154 13492 19654
rect 13740 19446 13768 19926
rect 13832 19553 13860 22063
rect 13924 21078 13952 22102
rect 14096 21956 14148 21962
rect 14096 21898 14148 21904
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13924 20806 13952 21014
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14016 20534 14044 21422
rect 14108 21010 14136 21898
rect 14200 21457 14228 22374
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14292 21690 14320 21830
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14186 21448 14242 21457
rect 14186 21383 14242 21392
rect 14200 21049 14228 21383
rect 14186 21040 14242 21049
rect 14096 21004 14148 21010
rect 14292 21010 14320 21626
rect 14186 20975 14242 20984
rect 14280 21004 14332 21010
rect 14096 20946 14148 20952
rect 14280 20946 14332 20952
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14108 20058 14136 20334
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14108 19854 14136 19994
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13818 19544 13874 19553
rect 14016 19514 14044 19654
rect 13818 19479 13874 19488
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 14292 19378 14320 20470
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 12990 18119 13046 18128
rect 12808 18090 12860 18096
rect 12820 18057 12848 18090
rect 12806 18048 12862 18057
rect 12806 17983 12862 17992
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17270 13400 18142
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 12900 17128 12952 17134
rect 12820 17076 12900 17082
rect 12820 17070 12952 17076
rect 12820 17054 12940 17070
rect 12820 16028 12848 17054
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13280 16114 13308 16594
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12992 16040 13044 16046
rect 12820 16000 12992 16028
rect 12992 15982 13044 15988
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13280 15094 13308 15438
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 14657 12848 14962
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12806 14648 12862 14657
rect 12950 14651 13258 14660
rect 12806 14583 12862 14592
rect 13372 14498 13400 17206
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16658 13492 16934
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 15706 13492 16594
rect 13556 16522 13584 19110
rect 13740 18970 13768 19110
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13832 18465 13860 19314
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13910 19000 13966 19009
rect 13910 18935 13966 18944
rect 13818 18456 13874 18465
rect 13818 18391 13874 18400
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17882 13860 18022
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13924 17762 13952 18935
rect 14016 18358 14044 19246
rect 14108 18601 14136 19246
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 14094 18592 14150 18601
rect 14094 18527 14150 18536
rect 14200 18426 14228 19178
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14016 17814 14044 18294
rect 13832 17734 13952 17762
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 16658 13676 17614
rect 13832 17610 13860 17734
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13912 17604 13964 17610
rect 13912 17546 13964 17552
rect 13726 17232 13782 17241
rect 13726 17167 13782 17176
rect 13740 17066 13768 17167
rect 13728 17060 13780 17066
rect 13728 17002 13780 17008
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13832 16561 13860 16934
rect 13818 16552 13874 16561
rect 13544 16516 13596 16522
rect 13818 16487 13874 16496
rect 13544 16458 13596 16464
rect 13634 16416 13690 16425
rect 13634 16351 13690 16360
rect 13648 15978 13676 16351
rect 13818 16280 13874 16289
rect 13818 16215 13874 16224
rect 13832 16182 13860 16215
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13832 15910 13860 16118
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13544 15360 13596 15366
rect 13542 15328 13544 15337
rect 13596 15328 13598 15337
rect 13542 15263 13598 15272
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14822 13584 14962
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13280 14470 13400 14498
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 12714 14376 12770 14385
rect 12714 14311 12770 14320
rect 13280 14074 13308 14470
rect 13358 14104 13414 14113
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13268 14068 13320 14074
rect 13358 14039 13360 14048
rect 13268 14010 13320 14016
rect 13412 14039 13414 14048
rect 13360 14010 13412 14016
rect 12912 13870 12940 14010
rect 13556 14006 13584 14486
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 12900 13864 12952 13870
rect 12898 13832 12900 13841
rect 12952 13832 12954 13841
rect 12716 13796 12768 13802
rect 12898 13767 12954 13776
rect 12716 13738 12768 13744
rect 12728 13308 12756 13738
rect 12806 13696 12862 13705
rect 12806 13631 12862 13640
rect 12820 13376 12848 13631
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13358 13560 13414 13569
rect 13358 13495 13414 13504
rect 13372 13444 13400 13495
rect 13648 13462 13676 15506
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 14618 13768 14894
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13728 14340 13780 14346
rect 13832 14328 13860 15846
rect 13924 15201 13952 17546
rect 14292 17542 14320 18634
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14108 17202 14136 17478
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 13910 15192 13966 15201
rect 13910 15127 13966 15136
rect 13910 14920 13966 14929
rect 13910 14855 13912 14864
rect 13964 14855 13966 14864
rect 13912 14826 13964 14832
rect 13780 14300 13860 14328
rect 13728 14282 13780 14288
rect 13740 13870 13768 14282
rect 13910 14240 13966 14249
rect 13910 14175 13966 14184
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13280 13416 13400 13444
rect 13636 13456 13688 13462
rect 12820 13348 13032 13376
rect 12728 13280 12848 13308
rect 12714 13016 12770 13025
rect 12714 12951 12716 12960
rect 12768 12951 12770 12960
rect 12716 12922 12768 12928
rect 12820 12782 12848 13280
rect 13004 12889 13032 13348
rect 12990 12880 13046 12889
rect 12990 12815 13046 12824
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 13280 12730 13308 13416
rect 13636 13398 13688 13404
rect 13358 13016 13414 13025
rect 13358 12951 13414 12960
rect 13542 13016 13598 13025
rect 13542 12951 13598 12960
rect 13372 12850 13400 12951
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13280 12702 13400 12730
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12728 11393 12756 12582
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12434 13400 12702
rect 13188 12406 13400 12434
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12714 11384 12770 11393
rect 12714 11319 12770 11328
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12636 10470 12664 11018
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12728 10146 12756 10678
rect 12636 10118 12756 10146
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12544 8265 12572 8502
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12360 7206 12388 7346
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12360 7041 12388 7142
rect 12346 7032 12402 7041
rect 12346 6967 12402 6976
rect 12636 6798 12664 10118
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 8974 12756 9862
rect 12820 9042 12848 12038
rect 13188 11665 13216 12406
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11354 13400 12038
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13464 11200 13492 11766
rect 13556 11393 13584 12951
rect 13542 11384 13598 11393
rect 13542 11319 13598 11328
rect 13372 11172 13492 11200
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12912 10742 12940 11086
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10810 13308 10950
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12912 10470 12940 10678
rect 13188 10470 13216 10746
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13268 9920 13320 9926
rect 13266 9888 13268 9897
rect 13320 9888 13322 9897
rect 13266 9823 13322 9832
rect 13266 9616 13322 9625
rect 13266 9551 13268 9560
rect 13320 9551 13322 9560
rect 13268 9522 13320 9528
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13372 9178 13400 11172
rect 13648 11098 13676 13398
rect 13740 13258 13768 13806
rect 13832 13802 13860 13942
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 12646 13768 13194
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13740 11354 13768 11834
rect 13832 11694 13860 12106
rect 13924 12102 13952 14175
rect 14016 13190 14044 16934
rect 14108 16697 14136 17138
rect 14200 16794 14228 17206
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14094 16688 14150 16697
rect 14094 16623 14150 16632
rect 14108 16182 14136 16623
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14096 16040 14148 16046
rect 14094 16008 14096 16017
rect 14148 16008 14150 16017
rect 14094 15943 14150 15952
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14094 15192 14150 15201
rect 14094 15127 14150 15136
rect 14108 15026 14136 15127
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14618 14136 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14200 14482 14228 15302
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14094 13152 14150 13161
rect 14094 13087 14150 13096
rect 14108 12374 14136 13087
rect 14186 12608 14242 12617
rect 14186 12543 14242 12552
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13912 12096 13964 12102
rect 14016 12073 14044 12310
rect 14096 12096 14148 12102
rect 13912 12038 13964 12044
rect 14002 12064 14058 12073
rect 14096 12038 14148 12044
rect 14002 11999 14058 12008
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14108 11608 14136 12038
rect 14016 11580 14136 11608
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13832 11218 13860 11494
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13464 11070 13676 11098
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13174 9072 13230 9081
rect 12808 9036 12860 9042
rect 13174 9007 13176 9016
rect 12808 8978 12860 8984
rect 13228 9007 13230 9016
rect 13360 9036 13412 9042
rect 13176 8978 13228 8984
rect 13360 8978 13412 8984
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12728 8378 12756 8910
rect 12806 8664 12862 8673
rect 12806 8599 12808 8608
rect 12860 8599 12862 8608
rect 12808 8570 12860 8576
rect 12728 8350 12848 8378
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 7954 12756 8230
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12360 6322 12388 6666
rect 12820 6322 12848 8350
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 7410 13400 8978
rect 13464 7886 13492 11070
rect 13634 10976 13690 10985
rect 13634 10911 13690 10920
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13556 10266 13584 10474
rect 13648 10266 13676 10911
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9654 13676 9862
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13360 7200 13412 7206
rect 13358 7168 13360 7177
rect 13412 7168 13414 7177
rect 12950 7100 13258 7109
rect 13358 7103 13414 7112
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 11980 6248 12032 6254
rect 13556 6225 13584 8366
rect 13648 8090 13676 8774
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13740 7546 13768 10542
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13832 7410 13860 11154
rect 13924 10849 13952 11494
rect 13910 10840 13966 10849
rect 13910 10775 13966 10784
rect 13924 9042 13952 10775
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13924 8265 13952 8298
rect 13910 8256 13966 8265
rect 13910 8191 13966 8200
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 11980 6190 12032 6196
rect 13542 6216 13598 6225
rect 14016 6186 14044 11580
rect 14200 11506 14228 12543
rect 14108 11478 14228 11506
rect 14108 6662 14136 11478
rect 14186 11384 14242 11393
rect 14186 11319 14188 11328
rect 14240 11319 14242 11328
rect 14188 11290 14240 11296
rect 14292 9722 14320 17138
rect 14384 16658 14412 23598
rect 14476 23225 14504 24142
rect 14554 24103 14610 24112
rect 14462 23216 14518 23225
rect 14462 23151 14518 23160
rect 14568 23118 14596 24103
rect 14752 23730 14780 24210
rect 14844 24206 14872 24783
rect 15028 24750 15056 25978
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14844 23769 14872 24142
rect 14830 23760 14886 23769
rect 14740 23724 14792 23730
rect 14830 23695 14886 23704
rect 14740 23666 14792 23672
rect 14936 23338 14964 24618
rect 15028 23730 15056 24686
rect 15016 23724 15068 23730
rect 15016 23666 15068 23672
rect 14936 23310 15056 23338
rect 14556 23112 14608 23118
rect 14556 23054 14608 23060
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22438 14596 22918
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14568 22166 14596 22374
rect 14556 22160 14608 22166
rect 14556 22102 14608 22108
rect 14568 21554 14596 22102
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14568 20534 14596 21490
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14568 20058 14596 20470
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14464 18964 14516 18970
rect 14568 18952 14596 19994
rect 14516 18924 14596 18952
rect 14464 18906 14516 18912
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14476 17785 14504 17818
rect 14462 17776 14518 17785
rect 14568 17746 14596 18158
rect 14462 17711 14518 17720
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14476 16794 14504 17478
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14462 16416 14518 16425
rect 14462 16351 14518 16360
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14384 13802 14412 16118
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12102 14412 12582
rect 14476 12434 14504 16351
rect 14568 15026 14596 17682
rect 14660 17649 14688 21830
rect 14844 20942 14872 22714
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14936 21894 14964 22578
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14924 21616 14976 21622
rect 14924 21558 14976 21564
rect 14936 21010 14964 21558
rect 15028 21010 15056 23310
rect 15120 22166 15148 26200
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 15566 26143 15622 26152
rect 15292 24880 15344 24886
rect 15292 24822 15344 24828
rect 15304 23497 15332 24822
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 15396 24070 15424 24686
rect 15384 24064 15436 24070
rect 15384 24006 15436 24012
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 23866 15516 24006
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15290 23488 15346 23497
rect 15290 23423 15346 23432
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15580 22030 15608 26143
rect 15764 23798 15792 26200
rect 16026 24440 16082 24449
rect 16026 24375 16082 24384
rect 16040 24138 16068 24375
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15658 23488 15714 23497
rect 15658 23423 15714 23432
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14832 20936 14884 20942
rect 14738 20904 14794 20913
rect 14832 20878 14884 20884
rect 14738 20839 14794 20848
rect 14752 20806 14780 20839
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14752 18222 14780 19314
rect 14830 18864 14886 18873
rect 14830 18799 14886 18808
rect 14740 18216 14792 18222
rect 14740 18158 14792 18164
rect 14752 18086 14780 18158
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14844 17882 14872 18799
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14646 17640 14702 17649
rect 14646 17575 14702 17584
rect 14844 17202 14872 17818
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14936 17082 14964 20946
rect 15120 20641 15148 21830
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15106 20632 15162 20641
rect 15580 20602 15608 21286
rect 15672 21010 15700 23423
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 17038 26200 17094 27000
rect 17682 26330 17738 27000
rect 17328 26302 17738 26330
rect 16762 25936 16818 25945
rect 16762 25871 16818 25880
rect 16578 25664 16634 25673
rect 16578 25599 16634 25608
rect 16672 25628 16724 25634
rect 16212 24132 16264 24138
rect 16212 24074 16264 24080
rect 16224 23322 16252 24074
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16316 22982 16344 23598
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 21146 16068 21422
rect 16132 21146 16160 21830
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 16316 20942 16344 22170
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 15106 20567 15162 20576
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16040 20369 16068 20402
rect 16026 20360 16082 20369
rect 16026 20295 16082 20304
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15028 19786 15056 19994
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 15016 19440 15068 19446
rect 15016 19382 15068 19388
rect 15028 19174 15056 19382
rect 15212 19258 15240 20198
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15120 19230 15240 19258
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15016 18828 15068 18834
rect 15120 18816 15148 19230
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15068 18788 15148 18816
rect 15016 18770 15068 18776
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14752 17054 14964 17082
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14660 16522 14688 16730
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14660 16114 14688 16458
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14752 14906 14780 17054
rect 15028 16590 15056 18362
rect 15212 17814 15240 19110
rect 15474 18864 15530 18873
rect 15474 18799 15530 18808
rect 15488 18698 15516 18799
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14830 15736 14886 15745
rect 14830 15671 14886 15680
rect 14844 15570 14872 15671
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15028 15337 15056 16390
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15014 15328 15070 15337
rect 15014 15263 15070 15272
rect 14568 14878 14780 14906
rect 14568 12617 14596 14878
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13394 14688 14350
rect 15120 13546 15148 15982
rect 15212 15434 15240 17750
rect 15580 17270 15608 19994
rect 15750 19952 15806 19961
rect 15750 19887 15806 19896
rect 15764 19378 15792 19887
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15672 19145 15700 19314
rect 15658 19136 15714 19145
rect 15658 19071 15714 19080
rect 15934 18592 15990 18601
rect 15934 18527 15990 18536
rect 15948 18222 15976 18527
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15856 17678 15884 17818
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15750 17368 15806 17377
rect 15750 17303 15806 17312
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15028 13530 15148 13546
rect 15028 13524 15160 13530
rect 15028 13518 15108 13524
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14554 12608 14610 12617
rect 14554 12543 14610 12552
rect 14830 12608 14886 12617
rect 14830 12543 14886 12552
rect 14740 12436 14792 12442
rect 14476 12406 14688 12434
rect 14660 12345 14688 12406
rect 14740 12378 14792 12384
rect 14646 12336 14702 12345
rect 14646 12271 14702 12280
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14384 11812 14412 12038
rect 14464 11824 14516 11830
rect 14384 11784 14464 11812
rect 14384 11150 14412 11784
rect 14464 11766 14516 11772
rect 14660 11370 14688 12271
rect 14752 12238 14780 12378
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11762 14780 12174
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14476 11342 14688 11370
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14476 10826 14504 11342
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14384 10798 14504 10826
rect 14384 10198 14412 10798
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14186 9616 14242 9625
rect 14186 9551 14242 9560
rect 14200 9518 14228 9551
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 8906 14228 9318
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14372 8628 14424 8634
rect 14476 8616 14504 10678
rect 14660 10130 14688 11154
rect 14844 10810 14872 12543
rect 14936 12434 14964 12718
rect 15028 12594 15056 13518
rect 15108 13466 15160 13472
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12730 15148 13330
rect 15212 12986 15240 14311
rect 15304 14074 15332 16050
rect 15396 14482 15424 16934
rect 15672 16658 15700 17138
rect 15764 17082 15792 17303
rect 15856 17270 15884 17478
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15936 17128 15988 17134
rect 15764 17054 15884 17082
rect 15936 17070 15988 17076
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 15706 15516 16390
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15672 15570 15700 15914
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15120 12702 15240 12730
rect 15028 12566 15148 12594
rect 14936 12406 15056 12434
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10124 14700 10130
rect 14568 10084 14648 10112
rect 14568 9586 14596 10084
rect 14648 10066 14700 10072
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14424 8588 14504 8616
rect 14372 8570 14424 8576
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14200 7886 14228 8434
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14292 6798 14320 8434
rect 14752 8090 14780 10610
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 8090 14872 9454
rect 14936 8430 14964 10066
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14660 6458 14688 7686
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 13542 6151 13598 6160
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 3194 11100 4558
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13740 3738 13768 5714
rect 14568 5642 14596 5714
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 12452 3126 12480 3674
rect 13832 3126 13860 4490
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3126 14136 4014
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 10140 3052 10192 3058
rect 10060 3012 10140 3040
rect 8392 2994 8444 3000
rect 10140 2994 10192 3000
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9416 800 9444 2450
rect 9784 2446 9812 2926
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 11900 2378 11928 2790
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 12084 800 12112 2450
rect 12452 2446 12480 2790
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 14752 800 14780 5714
rect 15028 2582 15056 12406
rect 15120 9654 15148 12566
rect 15212 12306 15240 12702
rect 15396 12442 15424 13806
rect 15580 12986 15608 15438
rect 15658 14104 15714 14113
rect 15658 14039 15714 14048
rect 15672 13938 15700 14039
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13462 15700 13670
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15382 12064 15438 12073
rect 15382 11999 15438 12008
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11082 15240 11494
rect 15200 11076 15252 11082
rect 15252 11036 15332 11064
rect 15200 11018 15252 11024
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 7478 15148 8774
rect 15212 7546 15240 9930
rect 15304 7818 15332 11036
rect 15396 9518 15424 11999
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15396 7410 15424 9454
rect 15488 8673 15516 12786
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15580 9926 15608 11018
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9654 15608 9862
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15580 9110 15608 9590
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15474 8664 15530 8673
rect 15474 8599 15530 8608
rect 15580 8430 15608 9046
rect 15672 8498 15700 11290
rect 15764 10810 15792 16458
rect 15856 12434 15884 17054
rect 15948 15706 15976 17070
rect 16040 16969 16068 20295
rect 16212 19236 16264 19242
rect 16212 19178 16264 19184
rect 16224 18834 16252 19178
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16026 16960 16082 16969
rect 16026 16895 16082 16904
rect 16040 16114 16068 16895
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 13870 15976 14214
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 16040 13326 16068 15846
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12714 15976 13126
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 16132 12434 16160 18022
rect 16224 17746 16252 18770
rect 16304 18080 16356 18086
rect 16302 18048 16304 18057
rect 16356 18048 16358 18057
rect 16302 17983 16358 17992
rect 16408 17785 16436 20742
rect 16500 20097 16528 20946
rect 16486 20088 16542 20097
rect 16486 20023 16542 20032
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16500 19174 16528 19654
rect 16592 19378 16620 25599
rect 16672 25570 16724 25576
rect 16684 24886 16712 25570
rect 16776 25537 16804 25871
rect 16762 25528 16818 25537
rect 16762 25463 16818 25472
rect 16672 24880 16724 24886
rect 16672 24822 16724 24828
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16854 22944 16910 22953
rect 16854 22879 16910 22888
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16684 20602 16712 21490
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16394 17776 16450 17785
rect 16212 17740 16264 17746
rect 16394 17711 16450 17720
rect 16212 17682 16264 17688
rect 16500 17610 16528 18634
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16592 17082 16620 19314
rect 16684 17354 16712 19722
rect 16776 18902 16804 22442
rect 16868 19174 16896 22879
rect 16960 21486 16988 23666
rect 16948 21480 17000 21486
rect 16946 21448 16948 21457
rect 17000 21448 17002 21457
rect 16946 21383 17002 21392
rect 17052 21010 17080 26200
rect 17222 24848 17278 24857
rect 17222 24783 17278 24792
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 17144 23118 17172 24210
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 22438 17172 23054
rect 17236 22710 17264 24783
rect 17328 23050 17356 26302
rect 17682 26200 17738 26302
rect 17958 26344 18014 26353
rect 17958 26279 18014 26288
rect 17868 26104 17920 26110
rect 17868 26046 17920 26052
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17420 25022 17448 25842
rect 17408 25016 17460 25022
rect 17408 24958 17460 24964
rect 17420 23730 17448 24958
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17420 22817 17448 22986
rect 17406 22808 17462 22817
rect 17406 22743 17462 22752
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 17880 22234 17908 26046
rect 17972 25945 18000 26279
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19246 26480 19302 26489
rect 19246 26415 19302 26424
rect 17958 25936 18014 25945
rect 17958 25871 18014 25880
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17958 23216 18014 23225
rect 17958 23151 17960 23160
rect 18012 23151 18014 23160
rect 17960 23122 18012 23128
rect 18340 22982 18368 26200
rect 18878 24440 18934 24449
rect 18878 24375 18934 24384
rect 18892 24342 18920 24375
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18432 23050 18460 24074
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18432 22710 18460 22986
rect 18892 22778 18920 24278
rect 18984 23322 19012 26200
rect 19260 23798 19288 26415
rect 19614 26330 19670 27000
rect 19352 26302 19670 26330
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19076 23610 19104 23734
rect 19352 23610 19380 26302
rect 19614 26200 19670 26302
rect 20258 26330 20314 27000
rect 20258 26302 20576 26330
rect 20258 26200 20314 26302
rect 20074 24984 20130 24993
rect 20074 24919 20130 24928
rect 20088 24206 20116 24919
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19076 23582 19380 23610
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 19154 22944 19210 22953
rect 19154 22879 19210 22888
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 18432 22094 18460 22646
rect 18512 22432 18564 22438
rect 18972 22432 19024 22438
rect 18564 22380 18644 22386
rect 18512 22374 18644 22380
rect 18972 22374 19024 22380
rect 18524 22358 18644 22374
rect 17604 22066 18368 22094
rect 18432 22066 18552 22094
rect 17130 21720 17186 21729
rect 17130 21655 17186 21664
rect 17144 21486 17172 21655
rect 17132 21480 17184 21486
rect 17132 21422 17184 21428
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17500 21344 17552 21350
rect 17604 21321 17632 22066
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 17880 21570 17908 21898
rect 18340 21842 18368 22066
rect 18418 21856 18474 21865
rect 18340 21814 18418 21842
rect 17950 21788 18258 21797
rect 18418 21791 18474 21800
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17788 21554 17908 21570
rect 18524 21554 18552 22066
rect 17776 21548 17908 21554
rect 17828 21542 17908 21548
rect 18512 21548 18564 21554
rect 17776 21490 17828 21496
rect 18512 21490 18564 21496
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17684 21412 17736 21418
rect 17684 21354 17736 21360
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17500 21286 17552 21292
rect 17590 21312 17646 21321
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 17236 20874 17264 21286
rect 17420 21078 17448 21286
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16960 18834 16988 20538
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17052 19417 17080 20198
rect 17144 19990 17172 20198
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17038 19408 17094 19417
rect 17038 19343 17094 19352
rect 17144 18834 17172 19790
rect 17236 19310 17264 20810
rect 17512 20602 17540 21286
rect 17590 21247 17646 21256
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17696 20398 17724 21354
rect 17788 20534 17816 21354
rect 17880 21321 17908 21422
rect 17866 21312 17922 21321
rect 17866 21247 17922 21256
rect 18524 20942 18552 21490
rect 18616 21486 18644 22358
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18878 21992 18934 22001
rect 18800 21622 18828 21966
rect 18878 21927 18934 21936
rect 18892 21894 18920 21927
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17682 20224 17738 20233
rect 17682 20159 17738 20168
rect 17696 20058 17724 20159
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17328 19009 17356 19314
rect 17406 19272 17462 19281
rect 17406 19207 17462 19216
rect 17314 19000 17370 19009
rect 17314 18935 17370 18944
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 16948 18624 17000 18630
rect 16946 18592 16948 18601
rect 17000 18592 17002 18601
rect 16946 18527 17002 18536
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16854 18184 16910 18193
rect 16854 18119 16856 18128
rect 16908 18119 16910 18128
rect 16856 18090 16908 18096
rect 17052 17762 17080 18226
rect 16960 17734 17080 17762
rect 16684 17326 16896 17354
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16500 17054 16620 17082
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 15366 16252 16526
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 14958 16252 15302
rect 16316 15162 16344 16594
rect 16500 16250 16528 17054
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16316 14346 16344 14962
rect 16304 14340 16356 14346
rect 16304 14282 16356 14288
rect 16316 14006 16344 14282
rect 16408 14074 16436 15030
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16500 13802 16528 15846
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 15856 12406 16068 12434
rect 16132 12406 16252 12434
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15934 10568 15990 10577
rect 15934 10503 15936 10512
rect 15988 10503 15990 10512
rect 15936 10474 15988 10480
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 16040 7970 16068 12406
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 11354 16160 12174
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 8498 16160 10542
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15948 7942 16068 7970
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15948 6934 15976 7942
rect 16224 7886 16252 12406
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16316 11898 16344 11999
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16316 11218 16344 11630
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11286 16436 11494
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16316 10130 16344 10542
rect 16408 10198 16436 11222
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16500 8634 16528 12106
rect 16592 9058 16620 16934
rect 16684 13394 16712 17138
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 16969 16804 17002
rect 16762 16960 16818 16969
rect 16762 16895 16818 16904
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16868 16574 16896 17326
rect 16960 16726 16988 17734
rect 17236 17542 17264 18634
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17052 16574 17080 16934
rect 16868 16546 17080 16574
rect 16776 15570 16804 16526
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16868 15502 16896 16546
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16776 14890 16804 15370
rect 16868 15026 16896 15438
rect 17052 15162 17080 16186
rect 17144 15570 17172 17002
rect 17236 15881 17264 17478
rect 17328 16561 17356 18935
rect 17420 18630 17448 19207
rect 17776 18896 17828 18902
rect 17776 18838 17828 18844
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17406 18456 17462 18465
rect 17788 18426 17816 18838
rect 17406 18391 17462 18400
rect 17776 18420 17828 18426
rect 17314 16552 17370 16561
rect 17420 16538 17448 18391
rect 17880 18408 17908 20402
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18248 19990 18276 20198
rect 18236 19984 18288 19990
rect 17958 19952 18014 19961
rect 18236 19926 18288 19932
rect 17958 19887 17960 19896
rect 18012 19887 18014 19896
rect 17960 19858 18012 19864
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18340 19514 18368 19722
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18234 19408 18290 19417
rect 18234 19343 18236 19352
rect 18288 19343 18290 19352
rect 18236 19314 18288 19320
rect 18248 18630 18276 19314
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17880 18380 18368 18408
rect 17776 18362 17828 18368
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18248 17649 18276 18158
rect 18234 17640 18290 17649
rect 18234 17575 18290 17584
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17788 16590 17816 17070
rect 17776 16584 17828 16590
rect 17420 16510 17540 16538
rect 17776 16526 17828 16532
rect 17314 16487 17370 16496
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17316 15904 17368 15910
rect 17222 15872 17278 15881
rect 17316 15846 17368 15852
rect 17222 15807 17278 15816
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12782 16712 13194
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16672 11756 16724 11762
rect 16776 11744 16804 14826
rect 16960 14822 16988 14894
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16854 14512 16910 14521
rect 16854 14447 16910 14456
rect 16868 13462 16896 14447
rect 17052 14346 17080 15098
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17052 14006 17080 14282
rect 17144 14278 17172 15506
rect 17328 14618 17356 15846
rect 17420 15434 17448 16390
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17420 14464 17448 14894
rect 17328 14436 17448 14464
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17144 13938 17172 14214
rect 17222 14104 17278 14113
rect 17222 14039 17224 14048
rect 17276 14039 17278 14048
rect 17224 14010 17276 14016
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16868 11898 16896 13398
rect 17144 13394 17172 13874
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16960 11830 16988 13262
rect 17328 13190 17356 14436
rect 17512 13870 17540 16510
rect 17788 15706 17816 16526
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18248 14890 18276 15098
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17920 13960 18092 13988
rect 17868 13942 17920 13948
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17604 13790 18000 13818
rect 17604 13682 17632 13790
rect 17972 13734 18000 13790
rect 17512 13654 17632 13682
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17512 12986 17540 13654
rect 18064 13569 18092 13960
rect 18050 13560 18106 13569
rect 17592 13524 17644 13530
rect 18050 13495 18106 13504
rect 17592 13466 17644 13472
rect 17604 12986 17632 13466
rect 18064 13258 18092 13495
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18340 13190 18368 18380
rect 18432 18057 18460 20198
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18524 19514 18552 19654
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18616 19378 18644 21422
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20641 18828 20742
rect 18786 20632 18842 20641
rect 18786 20567 18842 20576
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18696 20256 18748 20262
rect 18694 20224 18696 20233
rect 18748 20224 18750 20233
rect 18694 20159 18750 20168
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 18766 18552 19110
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18616 18630 18644 18838
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18708 18630 18736 18770
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18418 18048 18474 18057
rect 18418 17983 18474 17992
rect 18524 16726 18552 18566
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18616 16658 18644 18158
rect 18694 16824 18750 16833
rect 18694 16759 18750 16768
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 14482 18460 16390
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18524 14618 18552 15914
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18418 13560 18474 13569
rect 18418 13495 18474 13504
rect 18432 13326 18460 13495
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17052 12170 17080 12718
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16724 11716 16804 11744
rect 16672 11698 16724 11704
rect 16684 10266 16712 11698
rect 17052 11694 17080 12106
rect 17040 11688 17092 11694
rect 16946 11656 17002 11665
rect 17040 11630 17092 11636
rect 16946 11591 17002 11600
rect 16960 10674 16988 11591
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9586 16896 10066
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16592 9030 16712 9058
rect 16868 9042 16896 9522
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16592 8634 16620 8842
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16040 7274 16068 7822
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16684 6118 16712 9030
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16776 8430 16804 8842
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16868 8294 16896 8366
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15120 4690 15148 5510
rect 16316 4826 16344 5578
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 16868 4146 16896 5850
rect 17052 5778 17080 11086
rect 17236 10742 17264 12242
rect 17512 11937 17540 12310
rect 17498 11928 17554 11937
rect 17498 11863 17554 11872
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 10130 17172 10610
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17236 9654 17264 10202
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17236 7970 17264 9590
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 8498 17356 9318
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17420 8090 17448 9930
rect 17604 8498 17632 12718
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17696 9058 17724 11630
rect 17788 9178 17816 13126
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18524 12850 18552 13738
rect 18616 13462 18644 15982
rect 18708 14618 18736 16759
rect 18800 15978 18828 20402
rect 18892 17513 18920 21422
rect 18984 20602 19012 22374
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 19168 20398 19196 22879
rect 19536 22710 19564 24074
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 20352 23656 20404 23662
rect 20352 23598 20404 23604
rect 19708 23520 19760 23526
rect 19800 23520 19852 23526
rect 19708 23462 19760 23468
rect 19798 23488 19800 23497
rect 19852 23488 19854 23497
rect 19720 23186 19748 23462
rect 19798 23423 19854 23432
rect 20364 23186 20392 23598
rect 20456 23186 20484 23734
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 19524 22704 19576 22710
rect 19524 22646 19576 22652
rect 19720 22642 19748 23122
rect 20456 22710 20484 23122
rect 19984 22704 20036 22710
rect 19982 22672 19984 22681
rect 20444 22704 20496 22710
rect 20036 22672 20038 22681
rect 19708 22636 19760 22642
rect 20444 22646 20496 22652
rect 19982 22607 20038 22616
rect 19708 22578 19760 22584
rect 19614 22264 19670 22273
rect 19340 22228 19392 22234
rect 19614 22199 19670 22208
rect 19340 22170 19392 22176
rect 19352 21894 19380 22170
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19260 21570 19288 21830
rect 19340 21616 19392 21622
rect 19260 21564 19340 21570
rect 19260 21558 19392 21564
rect 19260 21542 19380 21558
rect 19260 20942 19288 21542
rect 19444 21010 19472 22034
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19536 21729 19564 21898
rect 19628 21894 19656 22199
rect 19720 22098 19748 22578
rect 20456 22234 20484 22646
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20548 22098 20576 26302
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26330 22246 27000
rect 22112 26302 22246 26330
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 23050 20668 25094
rect 20916 24274 20944 26200
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21192 23730 21220 24686
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21376 23798 21404 24550
rect 21560 24274 21588 26200
rect 22008 25084 22060 25090
rect 22008 25026 22060 25032
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21822 24032 21878 24041
rect 21822 23967 21878 23976
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21836 23254 21864 23967
rect 21824 23248 21876 23254
rect 21824 23190 21876 23196
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 21468 22234 21496 22374
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21836 22166 21864 23190
rect 20628 22160 20680 22166
rect 20628 22102 20680 22108
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19522 21720 19578 21729
rect 19522 21655 19578 21664
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19628 20964 19840 20992
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19260 19514 19288 20878
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19260 19292 19288 19450
rect 19352 19446 19380 20946
rect 19628 20874 19656 20964
rect 19616 20868 19668 20874
rect 19812 20856 19840 20964
rect 19984 20868 20036 20874
rect 19812 20828 19984 20856
rect 19616 20810 19668 20816
rect 19984 20810 20036 20816
rect 19432 20800 19484 20806
rect 19430 20768 19432 20777
rect 19484 20768 19486 20777
rect 19430 20703 19486 20712
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19628 20233 19656 20402
rect 19706 20360 19762 20369
rect 19706 20295 19708 20304
rect 19760 20295 19762 20304
rect 19708 20266 19760 20272
rect 19614 20224 19670 20233
rect 19614 20159 19670 20168
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19260 19264 19380 19292
rect 19352 18970 19380 19264
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19260 18426 19288 18906
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18878 17504 18934 17513
rect 18878 17439 18934 17448
rect 18984 16794 19012 18158
rect 19444 18086 19472 19926
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19628 18306 19656 19858
rect 20088 19854 20116 21830
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20180 20233 20208 20946
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20166 20224 20222 20233
rect 20166 20159 20222 20168
rect 20180 19922 20208 20159
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19720 18766 19748 19246
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19812 18601 19840 19654
rect 19798 18592 19854 18601
rect 19798 18527 19854 18536
rect 19628 18278 19748 18306
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19340 18080 19392 18086
rect 19338 18048 19340 18057
rect 19432 18080 19484 18086
rect 19392 18048 19394 18057
rect 19432 18022 19484 18028
rect 19338 17983 19394 17992
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19260 17649 19288 17818
rect 19246 17640 19302 17649
rect 19246 17575 19302 17584
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18892 15450 18920 16662
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19076 16250 19104 16390
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18984 15706 19012 15914
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19076 15586 19104 16050
rect 19168 15745 19196 16594
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19154 15736 19210 15745
rect 19154 15671 19210 15680
rect 18800 15422 18920 15450
rect 18984 15558 19104 15586
rect 18984 15434 19012 15558
rect 18972 15428 19024 15434
rect 18800 14890 18828 15422
rect 18972 15370 19024 15376
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18248 12702 18460 12730
rect 18248 12646 18276 12702
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18248 12186 18276 12378
rect 18340 12306 18368 12582
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18248 12158 18368 12186
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11762 17908 12038
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10742 17908 11018
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17880 9994 17908 10678
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17696 9030 17816 9058
rect 17788 8838 17816 9030
rect 18340 8974 18368 12158
rect 18432 11286 18460 12702
rect 18708 12617 18736 14282
rect 18892 14074 18920 15302
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18984 13802 19012 15370
rect 19168 15337 19196 15671
rect 19260 15366 19288 16526
rect 19248 15360 19300 15366
rect 19154 15328 19210 15337
rect 19248 15302 19300 15308
rect 19154 15263 19210 15272
rect 19352 15094 19380 17983
rect 19444 17678 19472 18022
rect 19628 17678 19656 18090
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19628 17134 19656 17614
rect 19616 17128 19668 17134
rect 19720 17105 19748 18278
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19812 18057 19840 18158
rect 19798 18048 19854 18057
rect 19798 17983 19854 17992
rect 19616 17070 19668 17076
rect 19706 17096 19762 17105
rect 19706 17031 19762 17040
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19812 16522 19840 17002
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19444 15570 19472 16118
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18786 13560 18842 13569
rect 18786 13495 18842 13504
rect 18694 12608 18750 12617
rect 18694 12543 18750 12552
rect 18800 12442 18828 13495
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18984 11558 19012 12718
rect 19076 12374 19104 14214
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 11370 19012 11494
rect 18984 11342 19104 11370
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18880 10532 18932 10538
rect 18880 10474 18932 10480
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17144 7954 17264 7970
rect 17132 7948 17264 7954
rect 17184 7942 17264 7948
rect 17132 7890 17184 7896
rect 17788 7818 17816 8774
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18432 7886 18460 10406
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18708 9654 18736 9862
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18524 8265 18552 9522
rect 18708 8634 18736 9590
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18708 8430 18736 8570
rect 18892 8498 18920 10474
rect 18984 9518 19012 11222
rect 19076 10606 19104 11342
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 19168 9382 19196 14826
rect 19444 14822 19472 14962
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19352 14634 19380 14758
rect 19260 14618 19380 14634
rect 19248 14612 19380 14618
rect 19300 14606 19380 14612
rect 19248 14554 19300 14560
rect 19260 14074 19288 14554
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19352 12434 19380 14418
rect 19260 12406 19380 12434
rect 19260 11354 19288 12406
rect 19444 12356 19472 14758
rect 19536 12918 19564 15098
rect 19628 15094 19656 15846
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19720 13394 19748 14962
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19524 12912 19576 12918
rect 19904 12889 19932 19722
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19996 18698 20024 19246
rect 20088 18970 20116 19246
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20180 18834 20208 19858
rect 20364 19786 20392 20742
rect 20640 20058 20668 22102
rect 21086 21856 21142 21865
rect 21086 21791 21142 21800
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20732 21078 20760 21286
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20732 19786 20760 20470
rect 20352 19780 20404 19786
rect 20720 19780 20772 19786
rect 20352 19722 20404 19728
rect 20548 19740 20720 19768
rect 20350 19680 20406 19689
rect 20350 19615 20406 19624
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 15201 20024 18226
rect 20088 17678 20116 18294
rect 20166 18048 20222 18057
rect 20166 17983 20222 17992
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20180 17610 20208 17983
rect 20272 17898 20300 19382
rect 20364 18222 20392 19615
rect 20548 19446 20576 19740
rect 20640 19514 20668 19740
rect 20720 19722 20772 19728
rect 20824 19514 20852 21490
rect 20916 21457 20944 21490
rect 21100 21457 21128 21791
rect 20902 21448 20958 21457
rect 20902 21383 20958 21392
rect 21086 21448 21142 21457
rect 21086 21383 21142 21392
rect 21456 21344 21508 21350
rect 21178 21312 21234 21321
rect 21456 21286 21508 21292
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21178 21247 21234 21256
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21100 20369 21128 20742
rect 21086 20360 21142 20369
rect 20996 20324 21048 20330
rect 21086 20295 21142 20304
rect 20996 20266 21048 20272
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20536 19440 20588 19446
rect 20588 19388 20760 19394
rect 20536 19382 20760 19388
rect 20548 19366 20760 19382
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20364 18086 20392 18158
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20272 17870 20392 17898
rect 20258 17640 20314 17649
rect 20168 17604 20220 17610
rect 20258 17575 20260 17584
rect 20168 17546 20220 17552
rect 20312 17575 20314 17584
rect 20260 17546 20312 17552
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16794 20116 16934
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20180 15570 20208 15914
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19982 15192 20038 15201
rect 19982 15127 20038 15136
rect 19996 14618 20024 15127
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19996 14278 20024 14554
rect 20088 14385 20116 15302
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20074 14376 20130 14385
rect 20074 14311 20130 14320
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19524 12854 19576 12860
rect 19890 12880 19946 12889
rect 19352 12328 19472 12356
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19260 8634 19288 11154
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18510 8256 18566 8265
rect 18510 8191 18566 8200
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 17420 800 17448 4626
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18524 3058 18552 6598
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18616 4078 18644 5034
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 19352 3466 19380 12328
rect 19536 12306 19564 12854
rect 19890 12815 19946 12824
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11082 19472 12174
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 19536 11694 19564 12106
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 9178 19472 11018
rect 19536 10810 19564 11630
rect 19996 11354 20024 11630
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19536 10470 19564 10746
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10130 19564 10406
rect 20180 10266 20208 14418
rect 20272 14113 20300 17274
rect 20364 14385 20392 17870
rect 20456 17814 20484 18022
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20548 17202 20576 19366
rect 20732 19310 20760 19366
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20640 19156 20668 19246
rect 21008 19156 21036 20266
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 20640 19128 21036 19156
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20824 17746 20852 18566
rect 20904 18080 20956 18086
rect 21100 18057 21128 19654
rect 20904 18022 20956 18028
rect 21086 18048 21142 18057
rect 20916 17814 20944 18022
rect 21086 17983 21142 17992
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20444 16516 20496 16522
rect 20548 16504 20576 17138
rect 20640 16998 20668 17682
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20718 16960 20774 16969
rect 20718 16895 20774 16904
rect 20732 16726 20760 16895
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20496 16476 20576 16504
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20444 16458 20496 16464
rect 20548 16182 20576 16476
rect 20536 16176 20588 16182
rect 20588 16124 20668 16130
rect 20536 16118 20668 16124
rect 20444 16108 20496 16114
rect 20548 16102 20668 16118
rect 20444 16050 20496 16056
rect 20350 14376 20406 14385
rect 20350 14311 20406 14320
rect 20258 14104 20314 14113
rect 20456 14074 20484 16050
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20548 15638 20576 15982
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20640 15450 20668 16102
rect 20732 15910 20760 16487
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20548 15434 20668 15450
rect 20548 15428 20680 15434
rect 20548 15422 20628 15428
rect 20548 15094 20576 15422
rect 20628 15370 20680 15376
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20640 14618 20668 15098
rect 20732 14958 20760 15098
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20258 14039 20314 14048
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12918 20300 13262
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 20548 8906 20576 13874
rect 20640 12900 20668 14010
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20732 13530 20760 13942
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20720 12912 20772 12918
rect 20640 12872 20720 12900
rect 20720 12854 20772 12860
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11830 20760 12038
rect 20720 11824 20772 11830
rect 20824 11801 20852 17682
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20994 17096 21050 17105
rect 20994 17031 21050 17040
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16561 20944 16934
rect 20902 16552 20958 16561
rect 20902 16487 20958 16496
rect 21008 15688 21036 17031
rect 21100 16658 21128 17614
rect 21192 17218 21220 21247
rect 21468 18834 21496 21286
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21284 17338 21312 18158
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21376 17542 21404 18022
rect 21454 17912 21510 17921
rect 21454 17847 21510 17856
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21192 17190 21404 17218
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 20916 15660 21036 15688
rect 20916 14278 20944 15660
rect 21100 15570 21128 16594
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21008 14958 21036 15506
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14346 21036 14758
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21100 14328 21128 15370
rect 21192 14929 21220 17002
rect 21376 16946 21404 17190
rect 21468 17105 21496 17847
rect 21454 17096 21510 17105
rect 21454 17031 21510 17040
rect 21376 16918 21496 16946
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21284 15162 21312 16458
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 21376 15162 21404 15370
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21468 15042 21496 16918
rect 21560 16114 21588 21286
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 21836 20874 21864 21082
rect 21640 20868 21692 20874
rect 21640 20810 21692 20816
rect 21824 20868 21876 20874
rect 21824 20810 21876 20816
rect 21652 20777 21680 20810
rect 21638 20768 21694 20777
rect 21638 20703 21694 20712
rect 21914 20088 21970 20097
rect 21914 20023 21916 20032
rect 21968 20023 21970 20032
rect 21916 19994 21968 20000
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21730 19136 21786 19145
rect 21730 19071 21786 19080
rect 21744 17882 21772 19071
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21638 17640 21694 17649
rect 21638 17575 21640 17584
rect 21692 17575 21694 17584
rect 21640 17546 21692 17552
rect 21744 16998 21772 17818
rect 21836 17542 21864 18770
rect 21928 17882 21956 19246
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21928 17542 21956 17818
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21836 17270 21864 17478
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21836 16658 21864 17206
rect 21916 16992 21968 16998
rect 21916 16934 21968 16940
rect 21928 16658 21956 16934
rect 21824 16652 21876 16658
rect 21824 16594 21876 16600
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21836 16017 21864 16594
rect 21822 16008 21878 16017
rect 21822 15943 21878 15952
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15366 21772 15846
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21284 15014 21496 15042
rect 21178 14920 21234 14929
rect 21178 14855 21234 14864
rect 21180 14340 21232 14346
rect 21100 14300 21180 14328
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13870 20944 14214
rect 21008 14074 21036 14282
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20720 11766 20772 11772
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20640 10470 20668 11086
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 5642 19472 8366
rect 19536 8362 19564 8774
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19536 5914 19564 8298
rect 20640 7410 20668 10406
rect 20916 9654 20944 13330
rect 21100 13258 21128 14300
rect 21180 14282 21232 14288
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21100 12850 21128 13194
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21284 12434 21312 15014
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21376 14414 21404 14826
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21836 14346 21864 14554
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 12434 21496 12786
rect 21100 12406 21312 12434
rect 21376 12406 21496 12434
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 21100 7342 21128 12406
rect 21376 12102 21404 12406
rect 21836 12102 21864 13738
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21376 11830 21404 12038
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21652 11082 21680 11766
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21192 9178 21220 11018
rect 21652 10810 21680 11018
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21284 10062 21312 10678
rect 21836 10674 21864 12038
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21928 10577 21956 13262
rect 21914 10568 21970 10577
rect 21914 10503 21970 10512
rect 21272 10056 21324 10062
rect 21732 10056 21784 10062
rect 21324 10004 21404 10010
rect 21272 9998 21404 10004
rect 21732 9998 21784 10004
rect 21284 9982 21404 9998
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 9518 21312 9862
rect 21376 9722 21404 9982
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21284 8974 21312 9454
rect 21744 9110 21772 9998
rect 22020 9738 22048 25026
rect 22112 18850 22140 26302
rect 22190 26200 22246 26302
rect 22834 26602 22890 27000
rect 23110 26616 23166 26625
rect 22834 26574 23110 26602
rect 22834 26200 22890 26574
rect 23110 26551 23166 26560
rect 23478 26330 23534 27000
rect 24122 26330 24178 27000
rect 24766 26330 24822 27000
rect 25134 26344 25190 26353
rect 23478 26302 23980 26330
rect 23478 26200 23534 26302
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22296 23186 22324 23802
rect 22466 23624 22522 23633
rect 22466 23559 22522 23568
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22296 21146 22324 21354
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 18970 22232 19110
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22112 18822 22232 18850
rect 22204 16674 22232 18822
rect 22388 16946 22416 21354
rect 22480 21010 22508 23559
rect 22572 23050 22600 25162
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23386 24440 23442 24449
rect 23386 24375 23442 24384
rect 23400 24342 23428 24375
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22664 23662 22692 23802
rect 23572 23792 23624 23798
rect 23572 23734 23624 23740
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22664 21486 22692 21966
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 19922 22692 20198
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22756 19854 22784 22510
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22466 19544 22522 19553
rect 22466 19479 22468 19488
rect 22520 19479 22522 19488
rect 22468 19450 22520 19456
rect 22572 18850 22600 19790
rect 22848 19514 22876 23598
rect 23296 23588 23348 23594
rect 23296 23530 23348 23536
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23032 22574 23060 23258
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 23124 22506 23152 23258
rect 23308 23186 23336 23530
rect 23584 23186 23612 23734
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23308 22710 23336 23122
rect 23584 23050 23612 23122
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23296 22704 23348 22710
rect 23480 22704 23532 22710
rect 23348 22652 23428 22658
rect 23296 22646 23428 22652
rect 23480 22646 23532 22652
rect 23308 22630 23428 22646
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23202 21856 23258 21865
rect 23202 21791 23258 21800
rect 23216 21622 23244 21791
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20777 23336 22102
rect 23400 21978 23428 22630
rect 23492 22545 23520 22646
rect 23478 22536 23534 22545
rect 23478 22471 23534 22480
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23400 21950 23520 21978
rect 23492 21570 23520 21950
rect 23584 21622 23612 22374
rect 23676 22030 23704 24006
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23768 22692 23796 23122
rect 23848 23112 23900 23118
rect 23846 23080 23848 23089
rect 23900 23080 23902 23089
rect 23846 23015 23902 23024
rect 23848 22704 23900 22710
rect 23768 22664 23848 22692
rect 23848 22646 23900 22652
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23400 21554 23520 21570
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23388 21548 23520 21554
rect 23440 21542 23520 21548
rect 23388 21490 23440 21496
rect 23492 21468 23520 21542
rect 23492 21440 23612 21468
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23294 20768 23350 20777
rect 23294 20703 23350 20712
rect 23400 20534 23428 21286
rect 23584 20806 23612 21440
rect 23662 21176 23718 21185
rect 23662 21111 23718 21120
rect 23676 21010 23704 21111
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23768 20874 23796 22374
rect 23860 21604 23888 22646
rect 23952 22094 23980 26302
rect 24122 26302 24624 26330
rect 24122 26200 24178 26302
rect 24492 24676 24544 24682
rect 24492 24618 24544 24624
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 24410 24440 24550
rect 24504 24410 24532 24618
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24030 23080 24086 23089
rect 24030 23015 24086 23024
rect 24044 22982 24072 23015
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 24596 22094 24624 26302
rect 24766 26302 25084 26330
rect 24766 26200 24822 26302
rect 25056 25838 25084 26302
rect 25134 26279 25190 26288
rect 25044 25832 25096 25838
rect 25044 25774 25096 25780
rect 24860 24608 24912 24614
rect 25148 24562 25176 26279
rect 25410 26200 25466 27000
rect 26054 26200 26110 27000
rect 26698 26330 26754 27000
rect 27342 26330 27398 27000
rect 26698 26302 27108 26330
rect 26698 26200 26754 26302
rect 24860 24550 24912 24556
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24688 22681 24716 23190
rect 24674 22672 24730 22681
rect 24674 22607 24730 22616
rect 23952 22066 24256 22094
rect 24596 22066 24716 22094
rect 23940 21616 23992 21622
rect 23860 21576 23940 21604
rect 23940 21558 23992 21564
rect 23952 20874 23980 21558
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23940 20868 23992 20874
rect 23940 20810 23992 20816
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23570 20632 23626 20641
rect 23570 20567 23572 20576
rect 23624 20567 23626 20576
rect 23848 20596 23900 20602
rect 23572 20538 23624 20544
rect 23848 20538 23900 20544
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23388 20392 23440 20398
rect 23756 20392 23808 20398
rect 23570 20360 23626 20369
rect 23440 20340 23570 20346
rect 23388 20334 23570 20340
rect 23400 20318 23570 20334
rect 23756 20334 23808 20340
rect 23570 20295 23626 20304
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22940 19258 22968 19654
rect 22848 19230 22968 19258
rect 22572 18822 22784 18850
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 17542 22508 18702
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22388 16918 22600 16946
rect 22204 16646 22416 16674
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 15094 22140 15506
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22112 14482 22140 15030
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22204 13938 22232 16390
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13530 22140 13670
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22204 13394 22232 13874
rect 22296 13569 22324 16526
rect 22282 13560 22338 13569
rect 22282 13495 22338 13504
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22204 12918 22232 13330
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21928 9710 22048 9738
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 20732 5778 20760 6734
rect 21928 6390 21956 9710
rect 22112 9654 22140 10950
rect 22204 10266 22232 12242
rect 22296 11830 22324 12242
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22020 8566 22048 9522
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22388 7857 22416 16646
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22480 15638 22508 15982
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22572 15065 22600 16918
rect 22664 16454 22692 18362
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22756 15978 22784 18822
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22558 15056 22614 15065
rect 22468 15020 22520 15026
rect 22558 14991 22614 15000
rect 22468 14962 22520 14968
rect 22480 14346 22508 14962
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14346 22600 14758
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22480 13530 22508 14010
rect 22848 13954 22876 19230
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23216 18426 23244 18634
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17542 23336 18702
rect 23400 18426 23428 18906
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23032 16522 23060 16730
rect 23020 16516 23072 16522
rect 23020 16458 23072 16464
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23216 16046 23244 16390
rect 23308 16250 23336 16730
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22572 13926 22876 13954
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22572 12434 22600 13926
rect 22652 13796 22704 13802
rect 22652 13738 22704 13744
rect 22480 12406 22600 12434
rect 22480 11121 22508 12406
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22466 11112 22522 11121
rect 22466 11047 22522 11056
rect 22572 10810 22600 12106
rect 22664 11286 22692 13738
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 23308 13274 23336 15302
rect 23400 15026 23428 18362
rect 23676 18358 23704 19654
rect 23768 19446 23796 20334
rect 23860 19514 23888 20538
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 23940 19236 23992 19242
rect 23940 19178 23992 19184
rect 23952 18834 23980 19178
rect 24044 18834 24072 19314
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23664 18352 23716 18358
rect 23716 18300 23796 18306
rect 23664 18294 23796 18300
rect 23676 18278 23796 18294
rect 23768 18222 23796 18278
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23662 17232 23718 17241
rect 23492 16998 23520 17206
rect 23662 17167 23718 17176
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 16114 23612 16934
rect 23676 16454 23704 17167
rect 23768 16590 23796 17682
rect 23860 17610 23888 18566
rect 23938 18048 23994 18057
rect 23938 17983 23994 17992
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23952 17270 23980 17983
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 17270 24072 17818
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23940 17128 23992 17134
rect 24044 17105 24072 17206
rect 23940 17070 23992 17076
rect 24030 17096 24086 17105
rect 23952 16658 23980 17070
rect 24030 17031 24086 17040
rect 24136 16794 24164 17478
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15434 23612 15846
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23584 15178 23612 15370
rect 23676 15337 23704 15370
rect 23662 15328 23718 15337
rect 23662 15263 23718 15272
rect 23584 15150 23704 15178
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23676 14414 23704 15150
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23386 13560 23442 13569
rect 23386 13495 23388 13504
rect 23440 13495 23442 13504
rect 23388 13466 23440 13472
rect 23216 13246 23336 13274
rect 23216 12918 23244 13246
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23204 12912 23256 12918
rect 23204 12854 23256 12860
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 23296 12436 23348 12442
rect 23400 12434 23428 12582
rect 23348 12406 23428 12434
rect 23492 12434 23520 13874
rect 23676 13190 23704 14350
rect 23754 13560 23810 13569
rect 23754 13495 23810 13504
rect 23768 13394 23796 13495
rect 23860 13394 23888 15506
rect 23952 14414 23980 16594
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23952 13734 23980 14350
rect 24122 14104 24178 14113
rect 24122 14039 24124 14048
rect 24176 14039 24178 14048
rect 24124 14010 24176 14016
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23768 12434 23796 12854
rect 23492 12406 23612 12434
rect 23296 12378 23348 12384
rect 22756 11830 22784 12378
rect 23584 12374 23612 12406
rect 23676 12406 23796 12434
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 23676 12238 23704 12406
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23676 11830 23704 12174
rect 23860 12102 23888 13330
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 22744 11824 22796 11830
rect 22744 11766 22796 11772
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22652 11280 22704 11286
rect 22652 11222 22704 11228
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22664 10674 22692 11222
rect 23676 11082 23704 11766
rect 23952 11558 23980 13330
rect 24228 12753 24256 22066
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24320 20942 24348 21966
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24320 20806 24348 20878
rect 24308 20800 24360 20806
rect 24308 20742 24360 20748
rect 24320 20398 24348 20742
rect 24504 20534 24532 21830
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24308 20392 24360 20398
rect 24308 20334 24360 20340
rect 24320 19718 24348 20334
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24412 17626 24440 18226
rect 24320 17610 24440 17626
rect 24308 17604 24440 17610
rect 24360 17598 24440 17604
rect 24308 17546 24360 17552
rect 24308 15428 24360 15434
rect 24308 15370 24360 15376
rect 24320 14822 24348 15370
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24412 14822 24440 15302
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24320 13870 24348 14758
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24214 12744 24270 12753
rect 24214 12679 24270 12688
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22652 10124 22704 10130
rect 22652 10066 22704 10072
rect 22664 9654 22692 10066
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22374 7848 22430 7857
rect 22374 7783 22430 7792
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22572 6866 22600 7278
rect 22756 7177 22784 9658
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23676 8294 23704 11018
rect 23952 9586 23980 11494
rect 24044 11150 24072 12038
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24320 11014 24348 13398
rect 24412 13326 24440 14214
rect 24596 13938 24624 20742
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24492 13796 24544 13802
rect 24492 13738 24544 13744
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24504 13190 24532 13738
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24504 12434 24532 13126
rect 24688 13002 24716 22066
rect 24780 21706 24808 24006
rect 24872 22098 24900 24550
rect 25056 24534 25176 24562
rect 25056 24274 25084 24534
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 25148 23798 25176 24346
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25136 22976 25188 22982
rect 25134 22944 25136 22953
rect 25188 22944 25190 22953
rect 25134 22879 25190 22888
rect 25240 22574 25268 24210
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25332 23338 25360 24142
rect 25424 23497 25452 26200
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25410 23488 25466 23497
rect 25410 23423 25466 23432
rect 25332 23310 25452 23338
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25148 22098 25176 22170
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 24952 21888 25004 21894
rect 24950 21856 24952 21865
rect 25004 21856 25006 21865
rect 24950 21791 25006 21800
rect 24780 21690 25084 21706
rect 24780 21684 25096 21690
rect 24780 21678 25044 21684
rect 25044 21626 25096 21632
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20534 24900 20810
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24780 18154 24808 20198
rect 25056 19922 25084 21490
rect 25240 21321 25268 22510
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25332 21622 25360 22374
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25226 21312 25282 21321
rect 25226 21247 25282 21256
rect 25320 20392 25372 20398
rect 25424 20380 25452 23310
rect 25516 21962 25544 24754
rect 25870 24712 25926 24721
rect 25870 24647 25926 24656
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25700 23662 25728 24006
rect 25688 23656 25740 23662
rect 25688 23598 25740 23604
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25700 22506 25728 22918
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25792 22166 25820 22374
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25596 21956 25648 21962
rect 25596 21898 25648 21904
rect 25608 20806 25636 21898
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25372 20352 25452 20380
rect 25320 20334 25372 20340
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25056 18630 25084 19314
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 24768 18148 24820 18154
rect 24768 18090 24820 18096
rect 24766 17912 24822 17921
rect 24766 17847 24768 17856
rect 24820 17847 24822 17856
rect 24768 17818 24820 17824
rect 24872 17610 24900 18566
rect 25056 18426 25084 18566
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24964 17270 24992 17682
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24412 12406 24532 12434
rect 24596 12974 24716 13002
rect 24412 12102 24440 12406
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 11558 24440 12038
rect 24400 11552 24452 11558
rect 24400 11494 24452 11500
rect 24412 11082 24440 11494
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23676 7410 23704 8230
rect 24044 7546 24072 9522
rect 24320 9081 24348 10406
rect 24596 9722 24624 12974
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12170 24716 12582
rect 24780 12306 24808 16390
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24872 15094 24900 15982
rect 24964 15638 24992 16594
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24872 14550 24900 14758
rect 24860 14544 24912 14550
rect 24964 14521 24992 15574
rect 24860 14486 24912 14492
rect 24950 14512 25006 14521
rect 24872 14006 24900 14486
rect 24950 14447 25006 14456
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24964 13802 24992 14214
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13326 25084 13670
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25148 12434 25176 18566
rect 25240 16538 25268 19722
rect 25332 18086 25360 19858
rect 25792 19446 25820 19858
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25792 18834 25820 19382
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25884 17105 25912 24647
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25976 22982 26004 24006
rect 26068 23118 26096 26200
rect 26148 25084 26200 25090
rect 26148 25026 26200 25032
rect 26160 24206 26188 25026
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26330 24440 26386 24449
rect 26330 24375 26386 24384
rect 26344 24274 26372 24375
rect 26332 24268 26384 24274
rect 26332 24210 26384 24216
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26424 24200 26476 24206
rect 26424 24142 26476 24148
rect 26436 23526 26464 24142
rect 26620 23594 26648 24754
rect 26698 24712 26754 24721
rect 26698 24647 26754 24656
rect 26712 23769 26740 24647
rect 26882 24440 26938 24449
rect 26882 24375 26938 24384
rect 26792 24132 26844 24138
rect 26792 24074 26844 24080
rect 26804 23798 26832 24074
rect 26896 24041 26924 24375
rect 26976 24268 27028 24274
rect 26976 24210 27028 24216
rect 26988 24070 27016 24210
rect 26976 24064 27028 24070
rect 26882 24032 26938 24041
rect 26976 24006 27028 24012
rect 26882 23967 26938 23976
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 26792 23792 26844 23798
rect 26698 23760 26754 23769
rect 26988 23769 27016 23802
rect 26792 23734 26844 23740
rect 26974 23760 27030 23769
rect 26698 23695 26754 23704
rect 26974 23695 27030 23704
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26424 23520 26476 23526
rect 26424 23462 26476 23468
rect 26436 23186 26464 23462
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26068 21962 26096 22442
rect 26160 22409 26188 23054
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26344 22778 26372 22986
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 26146 22400 26202 22409
rect 26146 22335 26202 22344
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25976 21078 26004 21286
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25962 20088 26018 20097
rect 25962 20023 25964 20032
rect 26016 20023 26018 20032
rect 25964 19994 26016 20000
rect 26160 19786 26188 21626
rect 26252 20874 26280 21830
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26240 20256 26292 20262
rect 26344 20244 26372 22714
rect 26292 20216 26372 20244
rect 26240 20198 26292 20204
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26252 19553 26280 20198
rect 26436 20074 26464 22918
rect 26620 22522 26648 23530
rect 27080 23361 27108 26302
rect 27342 26302 27568 26330
rect 27342 26200 27398 26302
rect 27160 25016 27212 25022
rect 27160 24958 27212 24964
rect 27342 24984 27398 24993
rect 27066 23352 27122 23361
rect 27066 23287 27122 23296
rect 26528 22494 26648 22522
rect 26528 22438 26556 22494
rect 26516 22432 26568 22438
rect 26516 22374 26568 22380
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26528 20874 26556 21898
rect 26620 21865 26648 22374
rect 26606 21856 26662 21865
rect 26606 21791 26662 21800
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 26712 21010 26740 21354
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 21010 27016 21286
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26516 20868 26568 20874
rect 26516 20810 26568 20816
rect 26528 20534 26556 20810
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26436 20046 26740 20074
rect 26238 19544 26294 19553
rect 26238 19479 26240 19488
rect 26292 19479 26294 19488
rect 26332 19508 26384 19514
rect 26240 19450 26292 19456
rect 26332 19450 26384 19456
rect 26344 19281 26372 19450
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26330 19272 26386 19281
rect 26330 19207 26386 19216
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26240 19168 26292 19174
rect 26528 19122 26556 19314
rect 26292 19116 26556 19122
rect 26240 19110 26556 19116
rect 26160 18834 26188 19110
rect 26252 19094 26556 19110
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25976 18358 26004 18634
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 26252 18034 26280 19094
rect 26516 18080 26568 18086
rect 26252 18006 26372 18034
rect 26516 18022 26568 18028
rect 25870 17096 25926 17105
rect 25870 17031 25926 17040
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25240 16522 25360 16538
rect 25240 16516 25372 16522
rect 25240 16510 25320 16516
rect 25320 16458 25372 16464
rect 25700 15570 25728 16594
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 24964 12406 25176 12434
rect 24964 12374 24992 12406
rect 24952 12368 25004 12374
rect 24952 12310 25004 12316
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24952 12232 25004 12238
rect 25240 12186 25268 15302
rect 25608 15201 25636 15302
rect 25594 15192 25650 15201
rect 25594 15127 25650 15136
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25004 12180 25268 12186
rect 24952 12174 25268 12180
rect 24676 12164 24728 12170
rect 24964 12158 25268 12174
rect 24676 12106 24728 12112
rect 24688 10062 24716 12106
rect 25516 11801 25544 14010
rect 25608 14006 25636 15127
rect 25700 14618 25728 15506
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 25700 13326 25728 14554
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25792 13190 25820 15302
rect 25872 14816 25924 14822
rect 25924 14764 26004 14770
rect 25872 14758 26004 14764
rect 25884 14742 26004 14758
rect 25976 14346 26004 14742
rect 25964 14340 26016 14346
rect 25964 14282 26016 14288
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25502 11792 25558 11801
rect 25136 11756 25188 11762
rect 25502 11727 25558 11736
rect 25136 11698 25188 11704
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24306 9072 24362 9081
rect 24306 9007 24362 9016
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24780 7993 24808 8978
rect 24766 7984 24822 7993
rect 24766 7919 24822 7928
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 22742 7168 22798 7177
rect 22742 7103 22798 7112
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 20732 5030 20760 5714
rect 22296 5370 22324 6258
rect 24044 6186 24072 7482
rect 25148 7313 25176 11698
rect 25884 11694 25912 12582
rect 25976 12442 26004 14282
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 25976 11218 26004 12378
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 26068 9450 26096 16594
rect 26160 15978 26188 17002
rect 26344 15994 26372 18006
rect 26528 17882 26556 18022
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26436 16182 26464 16526
rect 26424 16176 26476 16182
rect 26424 16118 26476 16124
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 26252 15966 26372 15994
rect 26252 15473 26280 15966
rect 26238 15464 26294 15473
rect 26148 15428 26200 15434
rect 26238 15399 26294 15408
rect 26148 15370 26200 15376
rect 26160 14890 26188 15370
rect 26528 15026 26556 16050
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26160 14074 26188 14826
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26252 13802 26280 14758
rect 26332 14544 26384 14550
rect 26332 14486 26384 14492
rect 26344 14074 26372 14486
rect 26528 14278 26556 14962
rect 26620 14822 26648 15642
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 12850 26280 13738
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26436 12782 26464 13126
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 25134 7304 25190 7313
rect 25134 7239 25190 7248
rect 24032 6180 24084 6186
rect 24032 6122 24084 6128
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 23492 5370 23520 5714
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23584 5234 23612 6054
rect 26252 5914 26280 8774
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 26712 5778 26740 20046
rect 26896 19786 26924 20470
rect 26988 20330 27016 20470
rect 27172 20398 27200 24958
rect 27342 24919 27398 24928
rect 27252 24064 27304 24070
rect 27252 24006 27304 24012
rect 27264 23186 27292 24006
rect 27252 23180 27304 23186
rect 27252 23122 27304 23128
rect 27264 22778 27292 23122
rect 27356 23032 27384 24919
rect 27540 24750 27568 26302
rect 27986 26200 28042 27000
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26330 29974 27000
rect 29918 26302 30328 26330
rect 29918 26200 29974 26302
rect 28000 25265 28028 26200
rect 27986 25256 28042 25265
rect 27986 25191 28042 25200
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27528 24744 27580 24750
rect 27528 24686 27580 24692
rect 27448 23798 27476 24686
rect 27712 24608 27764 24614
rect 27712 24550 27764 24556
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27436 23044 27488 23050
rect 27356 23004 27436 23032
rect 27436 22986 27488 22992
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27252 22568 27304 22574
rect 27252 22510 27304 22516
rect 27264 21554 27292 22510
rect 27540 22094 27568 23462
rect 27632 22506 27660 24278
rect 27724 24070 27752 24550
rect 28092 24274 28120 24550
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27712 23792 27764 23798
rect 27816 23780 27844 24074
rect 28092 24070 28120 24210
rect 28080 24064 28132 24070
rect 28080 24006 28132 24012
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27896 23792 27948 23798
rect 27816 23752 27896 23780
rect 27712 23734 27764 23740
rect 27896 23734 27948 23740
rect 27724 23508 27752 23734
rect 27804 23520 27856 23526
rect 27724 23480 27804 23508
rect 27804 23462 27856 23468
rect 27712 22976 27764 22982
rect 27710 22944 27712 22953
rect 27764 22944 27766 22953
rect 27710 22879 27766 22888
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27620 22500 27672 22506
rect 27620 22442 27672 22448
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 22234 27844 22374
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 28368 22166 28396 24210
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28552 23254 28580 24074
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28644 22953 28672 26200
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28828 23866 28856 24006
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28736 23225 28764 23666
rect 28920 23338 28948 24890
rect 29000 24880 29052 24886
rect 29000 24822 29052 24828
rect 29012 24313 29040 24822
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 29104 24342 29132 24686
rect 29288 24614 29316 26200
rect 29458 24848 29514 24857
rect 29458 24783 29514 24792
rect 30104 24812 30156 24818
rect 29368 24676 29420 24682
rect 29368 24618 29420 24624
rect 29184 24608 29236 24614
rect 29184 24550 29236 24556
rect 29276 24608 29328 24614
rect 29276 24550 29328 24556
rect 29092 24336 29144 24342
rect 28998 24304 29054 24313
rect 29092 24278 29144 24284
rect 28998 24239 29054 24248
rect 29104 24206 29132 24278
rect 29092 24200 29144 24206
rect 29092 24142 29144 24148
rect 29000 24064 29052 24070
rect 29196 24041 29224 24550
rect 29288 24274 29316 24550
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 29000 24006 29052 24012
rect 29182 24032 29238 24041
rect 29012 23662 29040 24006
rect 29182 23967 29238 23976
rect 29380 23905 29408 24618
rect 29366 23896 29422 23905
rect 29366 23831 29422 23840
rect 29380 23662 29408 23831
rect 29000 23656 29052 23662
rect 29000 23598 29052 23604
rect 29368 23656 29420 23662
rect 29368 23598 29420 23604
rect 29276 23588 29328 23594
rect 29276 23530 29328 23536
rect 28828 23310 28948 23338
rect 28722 23216 28778 23225
rect 28722 23151 28778 23160
rect 28630 22944 28686 22953
rect 28630 22879 28686 22888
rect 28828 22794 28856 23310
rect 29092 23248 29144 23254
rect 29092 23190 29144 23196
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28644 22766 28856 22794
rect 28920 22778 28948 23122
rect 29104 23050 29132 23190
rect 29092 23044 29144 23050
rect 29092 22986 29144 22992
rect 28908 22772 28960 22778
rect 28356 22160 28408 22166
rect 28356 22102 28408 22108
rect 27540 22066 27660 22094
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 27356 21486 27384 21898
rect 27434 21720 27490 21729
rect 27434 21655 27490 21664
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27448 20602 27476 21655
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27540 21146 27568 21490
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27160 20392 27212 20398
rect 27160 20334 27212 20340
rect 26976 20324 27028 20330
rect 26976 20266 27028 20272
rect 27540 20262 27568 20402
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27632 19922 27660 22066
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27710 21856 27766 21865
rect 27710 21791 27766 21800
rect 27724 21554 27752 21791
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27816 21486 27844 21966
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28644 21690 28672 22766
rect 28908 22714 28960 22720
rect 28814 22672 28870 22681
rect 28814 22607 28870 22616
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28538 21584 28594 21593
rect 28356 21548 28408 21554
rect 28538 21519 28594 21528
rect 28356 21490 28408 21496
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27710 20904 27766 20913
rect 27710 20839 27766 20848
rect 27724 19922 27752 20839
rect 27816 20058 27844 21422
rect 28368 21060 28396 21490
rect 28552 21185 28580 21519
rect 28538 21176 28594 21185
rect 28538 21111 28594 21120
rect 28368 21032 28580 21060
rect 28552 20942 28580 21032
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28540 20936 28592 20942
rect 28828 20913 28856 22607
rect 28920 22234 28948 22714
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28920 21350 28948 22170
rect 29104 21894 29132 22986
rect 29184 22432 29236 22438
rect 29184 22374 29236 22380
rect 29196 21962 29224 22374
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 28920 21146 28948 21286
rect 28908 21140 28960 21146
rect 28908 21082 28960 21088
rect 29104 20942 29132 21286
rect 29092 20936 29144 20942
rect 28540 20878 28592 20884
rect 28814 20904 28870 20913
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 28356 20460 28408 20466
rect 28356 20402 28408 20408
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27896 20052 27948 20058
rect 27896 19994 27948 20000
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26896 19334 26924 19722
rect 27908 19700 27936 19994
rect 28000 19854 28028 20402
rect 28080 20324 28132 20330
rect 28080 20266 28132 20272
rect 28092 19854 28120 20266
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 27816 19689 27936 19700
rect 27802 19680 27936 19689
rect 27858 19672 27936 19680
rect 27802 19615 27858 19624
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27618 19544 27674 19553
rect 27950 19547 28258 19556
rect 27618 19479 27674 19488
rect 26804 19306 26924 19334
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 26804 18766 26832 19306
rect 26882 19136 26938 19145
rect 26882 19071 26938 19080
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26804 18290 26832 18702
rect 26896 18601 26924 19071
rect 27264 18834 27292 19314
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 26882 18592 26938 18601
rect 26882 18527 26938 18536
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26804 18086 26832 18226
rect 26792 18080 26844 18086
rect 26792 18022 26844 18028
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 26804 17610 26832 18022
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26804 17270 26832 17546
rect 26792 17264 26844 17270
rect 26792 17206 26844 17212
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16590 27292 17070
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 16250 27292 16390
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26896 15094 26924 15506
rect 27172 15502 27200 16050
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26884 15088 26936 15094
rect 26884 15030 26936 15036
rect 26988 14958 27016 15302
rect 27448 15162 27476 18022
rect 27632 17882 27660 19479
rect 28368 19378 28396 20402
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 18426 27752 18566
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27816 17898 27844 19314
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 28368 18358 28396 19314
rect 28460 18902 28488 20878
rect 29092 20878 29144 20884
rect 28814 20839 28870 20848
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 28828 19990 28856 20742
rect 28816 19984 28868 19990
rect 28816 19926 28868 19932
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28630 19000 28686 19009
rect 28736 18970 28764 19654
rect 28920 19446 28948 19926
rect 29104 19922 29132 20878
rect 29184 20800 29236 20806
rect 29184 20742 29236 20748
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 28908 19440 28960 19446
rect 28908 19382 28960 19388
rect 28814 19272 28870 19281
rect 28814 19207 28870 19216
rect 28828 18970 28856 19207
rect 28630 18935 28686 18944
rect 28724 18964 28776 18970
rect 28644 18902 28672 18935
rect 28724 18906 28776 18912
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28448 18896 28500 18902
rect 28448 18838 28500 18844
rect 28632 18896 28684 18902
rect 28632 18838 28684 18844
rect 28644 18766 28672 18838
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27724 17870 27844 17898
rect 27724 17610 27752 17870
rect 28092 17746 28120 18226
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28354 17776 28410 17785
rect 27804 17740 27856 17746
rect 27804 17682 27856 17688
rect 28080 17740 28132 17746
rect 28354 17711 28410 17720
rect 28538 17776 28594 17785
rect 28538 17711 28594 17720
rect 28724 17740 28776 17746
rect 28080 17682 28132 17688
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27816 17202 27844 17682
rect 28368 17513 28396 17711
rect 28354 17504 28410 17513
rect 27950 17436 28258 17445
rect 28354 17439 28410 17448
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 28552 17105 28580 17711
rect 28724 17682 28776 17688
rect 28538 17096 28594 17105
rect 28538 17031 28594 17040
rect 27528 16992 27580 16998
rect 27528 16934 27580 16940
rect 27540 16640 27568 16934
rect 28736 16658 28764 17682
rect 27804 16652 27856 16658
rect 27540 16612 27804 16640
rect 27540 16114 27568 16612
rect 27804 16594 27856 16600
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27632 15502 27660 15846
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27618 15192 27674 15201
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27436 15156 27488 15162
rect 27618 15127 27674 15136
rect 27436 15098 27488 15104
rect 26976 14952 27028 14958
rect 26976 14894 27028 14900
rect 27172 14618 27200 15098
rect 27448 15026 27476 15098
rect 27632 15026 27660 15127
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27448 14822 27476 14962
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27724 14074 27752 15846
rect 27816 15434 27844 16118
rect 28736 15706 28764 16594
rect 28920 16114 28948 17818
rect 29012 16697 29040 18906
rect 28998 16688 29054 16697
rect 28998 16623 29054 16632
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 15162 27844 15370
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 26882 13696 26938 13705
rect 26882 13631 26938 13640
rect 26896 13161 26924 13631
rect 26882 13152 26938 13161
rect 26882 13087 26938 13096
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27816 9654 27844 11018
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 9648 27856 9654
rect 27804 9590 27856 9596
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24780 5302 24808 5578
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19904 4486 19932 4626
rect 20916 4622 20944 5170
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21376 4622 21404 5034
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 23584 4554 23612 5170
rect 25504 5092 25556 5098
rect 25504 5034 25556 5040
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19904 3126 19932 4422
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20088 800 20116 4014
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22756 800 22784 2926
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 25516 2650 25544 5034
rect 26712 3602 26740 5714
rect 27528 5636 27580 5642
rect 27528 5578 27580 5584
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 27356 4826 27384 5102
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 26700 3596 26752 3602
rect 26700 3538 26752 3544
rect 27540 2650 27568 5578
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 28552 5302 28580 15642
rect 28724 8832 28776 8838
rect 28724 8774 28776 8780
rect 28736 6390 28764 8774
rect 28724 6384 28776 6390
rect 28724 6326 28776 6332
rect 27620 5296 27672 5302
rect 27620 5238 27672 5244
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 27632 3534 27660 5238
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 28736 2514 28764 6326
rect 29104 5302 29132 19858
rect 29196 19310 29224 20742
rect 29288 19922 29316 23530
rect 29472 22817 29500 24783
rect 30104 24754 30156 24760
rect 30116 24206 30144 24754
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 29458 22808 29514 22817
rect 29458 22743 29514 22752
rect 29368 22092 29420 22098
rect 29368 22034 29420 22040
rect 29380 21894 29408 22034
rect 29368 21888 29420 21894
rect 29368 21830 29420 21836
rect 29380 21622 29408 21830
rect 29368 21616 29420 21622
rect 29368 21558 29420 21564
rect 29380 20942 29408 21558
rect 29368 20936 29420 20942
rect 29368 20878 29420 20884
rect 29380 20534 29408 20878
rect 29368 20528 29420 20534
rect 29368 20470 29420 20476
rect 29276 19916 29328 19922
rect 29276 19858 29328 19864
rect 29380 19718 29408 20470
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29380 19446 29408 19654
rect 29368 19440 29420 19446
rect 29420 19400 29500 19428
rect 29368 19382 29420 19388
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29380 18426 29408 19246
rect 29472 18630 29500 19400
rect 29840 19310 29868 24142
rect 30300 23882 30328 26302
rect 30562 26200 30618 27000
rect 30930 26616 30986 26625
rect 30986 26574 31064 26602
rect 30930 26551 30986 26560
rect 30576 24342 30604 26200
rect 30932 26172 30984 26178
rect 30932 26114 30984 26120
rect 30564 24336 30616 24342
rect 30564 24278 30616 24284
rect 30300 23854 30420 23882
rect 30392 23798 30420 23854
rect 30196 23792 30248 23798
rect 30196 23734 30248 23740
rect 30380 23792 30432 23798
rect 30380 23734 30432 23740
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30012 23656 30064 23662
rect 30012 23598 30064 23604
rect 30024 23186 30052 23598
rect 30116 23322 30144 23666
rect 30208 23322 30236 23734
rect 30104 23316 30156 23322
rect 30104 23258 30156 23264
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30012 23180 30064 23186
rect 30012 23122 30064 23128
rect 30380 22976 30432 22982
rect 30380 22918 30432 22924
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 30104 22704 30156 22710
rect 30104 22646 30156 22652
rect 30116 22522 30144 22646
rect 30116 22494 30236 22522
rect 30392 22506 30420 22918
rect 30562 22536 30618 22545
rect 30208 22438 30236 22494
rect 30380 22500 30432 22506
rect 30562 22471 30618 22480
rect 30380 22442 30432 22448
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30116 22030 30144 22374
rect 30208 22094 30236 22374
rect 30576 22166 30604 22471
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 30668 22098 30696 22918
rect 30288 22094 30340 22098
rect 30208 22092 30340 22094
rect 30208 22066 30288 22092
rect 30288 22034 30340 22040
rect 30656 22092 30708 22098
rect 30656 22034 30708 22040
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30378 21992 30434 22001
rect 30378 21927 30434 21936
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30024 21690 30052 21830
rect 30012 21684 30064 21690
rect 30012 21626 30064 21632
rect 30300 21554 30328 21830
rect 30288 21548 30340 21554
rect 30288 21490 30340 21496
rect 30300 21162 30328 21490
rect 30392 21321 30420 21927
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30484 21486 30512 21830
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30378 21312 30434 21321
rect 30378 21247 30434 21256
rect 30300 21134 30420 21162
rect 30196 20936 30248 20942
rect 30196 20878 30248 20884
rect 30208 20398 30236 20878
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30392 20330 30420 21134
rect 30668 21078 30696 21626
rect 30760 21622 30788 23734
rect 30944 23730 30972 26114
rect 31036 23730 31064 26574
rect 31206 26200 31262 27000
rect 31850 26330 31906 27000
rect 32126 26480 32182 26489
rect 32126 26415 32182 26424
rect 31850 26302 32076 26330
rect 31850 26200 31906 26302
rect 31220 24750 31248 26200
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31576 24404 31628 24410
rect 31576 24346 31628 24352
rect 31116 24200 31168 24206
rect 31116 24142 31168 24148
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 31024 23724 31076 23730
rect 31024 23666 31076 23672
rect 31128 23526 31156 24142
rect 31390 23624 31446 23633
rect 31390 23559 31446 23568
rect 31404 23526 31432 23559
rect 31116 23520 31168 23526
rect 31116 23462 31168 23468
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31128 22574 31156 23462
rect 31588 22982 31616 24346
rect 31668 24268 31720 24274
rect 31668 24210 31720 24216
rect 31680 23594 31708 24210
rect 31850 24032 31906 24041
rect 31850 23967 31906 23976
rect 31668 23588 31720 23594
rect 31668 23530 31720 23536
rect 31864 23526 31892 23967
rect 31852 23520 31904 23526
rect 31852 23462 31904 23468
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31576 22976 31628 22982
rect 31576 22918 31628 22924
rect 31576 22772 31628 22778
rect 31576 22714 31628 22720
rect 31668 22772 31720 22778
rect 31668 22714 31720 22720
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31024 22568 31076 22574
rect 31024 22510 31076 22516
rect 31116 22568 31168 22574
rect 31116 22510 31168 22516
rect 30840 22500 30892 22506
rect 30840 22442 30892 22448
rect 30852 22137 30880 22442
rect 30838 22128 30894 22137
rect 31036 22098 31064 22510
rect 31220 22250 31248 22578
rect 31588 22574 31616 22714
rect 31680 22681 31708 22714
rect 31666 22672 31722 22681
rect 31666 22607 31722 22616
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31772 22438 31800 23054
rect 31864 22642 31892 23462
rect 32048 23118 32076 26302
rect 31944 23112 31996 23118
rect 31944 23054 31996 23060
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31760 22432 31812 22438
rect 31760 22374 31812 22380
rect 31128 22222 31248 22250
rect 31128 22166 31156 22222
rect 31116 22160 31168 22166
rect 31116 22102 31168 22108
rect 30838 22063 30894 22072
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 30748 21616 30800 21622
rect 30748 21558 30800 21564
rect 30840 21412 30892 21418
rect 30840 21354 30892 21360
rect 30656 21072 30708 21078
rect 30656 21014 30708 21020
rect 30852 20942 30880 21354
rect 31036 21350 31064 21626
rect 31024 21344 31076 21350
rect 31024 21286 31076 21292
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 30380 20324 30432 20330
rect 30380 20266 30432 20272
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29828 18828 29880 18834
rect 29828 18770 29880 18776
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29368 18420 29420 18426
rect 29368 18362 29420 18368
rect 29472 18290 29500 18566
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29472 18086 29500 18226
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 29472 17678 29500 18022
rect 29460 17672 29512 17678
rect 29460 17614 29512 17620
rect 29368 17536 29420 17542
rect 29368 17478 29420 17484
rect 29380 16522 29408 17478
rect 29472 17270 29500 17614
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 29564 15910 29592 16526
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29564 12209 29592 15846
rect 29656 15609 29684 18294
rect 29748 16726 29776 18566
rect 29840 18426 29868 18770
rect 29932 18698 29960 20198
rect 30392 19854 30420 20266
rect 30380 19848 30432 19854
rect 30380 19790 30432 19796
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 29828 18420 29880 18426
rect 29828 18362 29880 18368
rect 30024 17746 30052 18770
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 30104 18692 30156 18698
rect 30104 18634 30156 18640
rect 30116 18057 30144 18634
rect 30102 18048 30158 18057
rect 30102 17983 30158 17992
rect 30208 17921 30236 18702
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30300 18222 30328 18566
rect 30288 18216 30340 18222
rect 30288 18158 30340 18164
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30194 17912 30250 17921
rect 30194 17847 30250 17856
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30024 17134 30052 17682
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17241 30236 17478
rect 30300 17338 30328 18022
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30194 17232 30250 17241
rect 30194 17167 30250 17176
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29736 16720 29788 16726
rect 29736 16662 29788 16668
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 29642 15600 29698 15609
rect 29642 15535 29698 15544
rect 29550 12200 29606 12209
rect 29550 12135 29606 12144
rect 30024 11665 30052 16594
rect 30392 16153 30420 17750
rect 30668 16561 30696 19314
rect 31128 18290 31156 22102
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 31484 20800 31536 20806
rect 31484 20742 31536 20748
rect 31496 20602 31524 20742
rect 31772 20602 31800 21082
rect 31864 20602 31892 22578
rect 31956 22234 31984 23054
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 31944 22228 31996 22234
rect 31944 22170 31996 22176
rect 31942 21992 31998 22001
rect 31942 21927 31944 21936
rect 31996 21927 31998 21936
rect 31944 21898 31996 21904
rect 32048 21418 32076 22374
rect 32140 21894 32168 26415
rect 32494 26200 32550 27000
rect 33138 26330 33194 27000
rect 33598 26344 33654 26353
rect 33138 26302 33548 26330
rect 33138 26200 33194 26302
rect 32404 25288 32456 25294
rect 32404 25230 32456 25236
rect 32220 24676 32272 24682
rect 32220 24618 32272 24624
rect 32232 23730 32260 24618
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32220 23520 32272 23526
rect 32220 23462 32272 23468
rect 32128 21888 32180 21894
rect 32128 21830 32180 21836
rect 32232 21554 32260 23462
rect 32310 23080 32366 23089
rect 32310 23015 32366 23024
rect 32324 22642 32352 23015
rect 32312 22636 32364 22642
rect 32312 22578 32364 22584
rect 32310 21584 32366 21593
rect 32220 21548 32272 21554
rect 32310 21519 32312 21528
rect 32220 21490 32272 21496
rect 32364 21519 32366 21528
rect 32312 21490 32364 21496
rect 32036 21412 32088 21418
rect 32036 21354 32088 21360
rect 32220 21412 32272 21418
rect 32220 21354 32272 21360
rect 32048 21146 32076 21354
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31852 20596 31904 20602
rect 31852 20538 31904 20544
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31220 19514 31248 20334
rect 31666 20088 31722 20097
rect 31666 20023 31722 20032
rect 31300 19984 31352 19990
rect 31300 19926 31352 19932
rect 31312 19514 31340 19926
rect 31680 19922 31708 20023
rect 31484 19916 31536 19922
rect 31484 19858 31536 19864
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31300 19508 31352 19514
rect 31300 19450 31352 19456
rect 31220 18766 31248 19450
rect 31404 19446 31432 19722
rect 31392 19440 31444 19446
rect 31392 19382 31444 19388
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30852 17882 30880 18158
rect 31128 17882 31156 18226
rect 30840 17876 30892 17882
rect 31116 17876 31168 17882
rect 30840 17818 30892 17824
rect 31036 17836 31116 17864
rect 31036 17678 31064 17836
rect 31116 17818 31168 17824
rect 31300 17740 31352 17746
rect 31300 17682 31352 17688
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 31312 17270 31340 17682
rect 31300 17264 31352 17270
rect 31300 17206 31352 17212
rect 30654 16552 30710 16561
rect 30654 16487 30710 16496
rect 30378 16144 30434 16153
rect 30378 16079 30434 16088
rect 30380 15972 30432 15978
rect 30380 15914 30432 15920
rect 30392 13938 30420 15914
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30010 11656 30066 11665
rect 30010 11591 30066 11600
rect 31312 11150 31340 17206
rect 31496 16726 31524 19858
rect 31576 19712 31628 19718
rect 31576 19654 31628 19660
rect 31588 18873 31616 19654
rect 31772 19378 31800 20538
rect 31864 20330 31892 20538
rect 31852 20324 31904 20330
rect 31852 20266 31904 20272
rect 32036 20256 32088 20262
rect 32036 20198 32088 20204
rect 31852 19440 31904 19446
rect 31852 19382 31904 19388
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31574 18864 31630 18873
rect 31574 18799 31630 18808
rect 31760 18148 31812 18154
rect 31760 18090 31812 18096
rect 31484 16720 31536 16726
rect 31484 16662 31536 16668
rect 31772 13705 31800 18090
rect 31758 13696 31814 13705
rect 31758 13631 31814 13640
rect 31864 12434 31892 19382
rect 32048 17649 32076 20198
rect 32140 19145 32168 21286
rect 32126 19136 32182 19145
rect 32126 19071 32182 19080
rect 32128 18828 32180 18834
rect 32128 18770 32180 18776
rect 32140 18630 32168 18770
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 32034 17640 32090 17649
rect 32034 17575 32090 17584
rect 32232 13258 32260 21354
rect 32416 21078 32444 25230
rect 32508 22234 32536 26200
rect 33324 25492 33376 25498
rect 33324 25434 33376 25440
rect 32772 25220 32824 25226
rect 32772 25162 32824 25168
rect 32680 25152 32732 25158
rect 32680 25094 32732 25100
rect 32586 23488 32642 23497
rect 32586 23423 32642 23432
rect 32600 23186 32628 23423
rect 32588 23180 32640 23186
rect 32588 23122 32640 23128
rect 32496 22228 32548 22234
rect 32496 22170 32548 22176
rect 32692 22094 32720 25094
rect 32784 24070 32812 25162
rect 32862 24984 32918 24993
rect 32862 24919 32918 24928
rect 32876 24410 32904 24919
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32864 24404 32916 24410
rect 32864 24346 32916 24352
rect 33048 24268 33100 24274
rect 33048 24210 33100 24216
rect 32772 24064 32824 24070
rect 32772 24006 32824 24012
rect 32862 23896 32918 23905
rect 32862 23831 32864 23840
rect 32916 23831 32918 23840
rect 32864 23802 32916 23808
rect 33060 23769 33088 24210
rect 33046 23760 33102 23769
rect 33046 23695 33102 23704
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32772 23316 32824 23322
rect 32772 23258 32824 23264
rect 32784 22409 32812 23258
rect 32956 23112 33008 23118
rect 32956 23054 33008 23060
rect 32968 22982 32996 23054
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 33232 22772 33284 22778
rect 33232 22714 33284 22720
rect 33244 22438 33272 22714
rect 33232 22432 33284 22438
rect 32770 22400 32826 22409
rect 33232 22374 33284 22380
rect 32770 22335 32826 22344
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32772 22094 32824 22098
rect 32692 22092 32824 22094
rect 32692 22066 32772 22092
rect 32772 22034 32824 22040
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32404 21072 32456 21078
rect 32404 21014 32456 21020
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32324 20233 32352 20402
rect 32310 20224 32366 20233
rect 32310 20159 32366 20168
rect 32416 20074 32444 21014
rect 32680 20528 32732 20534
rect 32784 20505 32812 21490
rect 33244 21418 33272 21626
rect 33232 21412 33284 21418
rect 33232 21354 33284 21360
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32862 21040 32918 21049
rect 33336 21010 33364 25434
rect 33520 24138 33548 26302
rect 33598 26279 33654 26288
rect 33782 26330 33838 27000
rect 33782 26302 34284 26330
rect 33508 24132 33560 24138
rect 33508 24074 33560 24080
rect 33612 24018 33640 26279
rect 33782 26200 33838 26302
rect 33968 26104 34020 26110
rect 33968 26046 34020 26052
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33520 23990 33640 24018
rect 33520 22094 33548 23990
rect 33888 23594 33916 24142
rect 33876 23588 33928 23594
rect 33876 23530 33928 23536
rect 33784 23520 33836 23526
rect 33784 23462 33836 23468
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33598 22808 33654 22817
rect 33598 22743 33654 22752
rect 33612 22506 33640 22743
rect 33704 22710 33732 22918
rect 33692 22704 33744 22710
rect 33692 22646 33744 22652
rect 33796 22574 33824 23462
rect 33888 22778 33916 23530
rect 33876 22772 33928 22778
rect 33876 22714 33928 22720
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33520 22066 33640 22094
rect 33414 21720 33470 21729
rect 33414 21655 33416 21664
rect 33468 21655 33470 21664
rect 33416 21626 33468 21632
rect 32862 20975 32864 20984
rect 32916 20975 32918 20984
rect 33324 21004 33376 21010
rect 32864 20946 32916 20952
rect 33324 20946 33376 20952
rect 32876 20602 32904 20946
rect 32864 20596 32916 20602
rect 32864 20538 32916 20544
rect 32680 20470 32732 20476
rect 32770 20496 32826 20505
rect 32324 20046 32444 20074
rect 32324 19310 32352 20046
rect 32402 19952 32458 19961
rect 32402 19887 32458 19896
rect 32416 19446 32444 19887
rect 32404 19440 32456 19446
rect 32404 19382 32456 19388
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 32404 19304 32456 19310
rect 32404 19246 32456 19252
rect 32416 18902 32444 19246
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32404 18896 32456 18902
rect 32404 18838 32456 18844
rect 32508 17814 32536 19110
rect 32588 18896 32640 18902
rect 32588 18838 32640 18844
rect 32496 17808 32548 17814
rect 32496 17750 32548 17756
rect 32600 16017 32628 18838
rect 32692 17513 32720 20470
rect 32770 20431 32826 20440
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33612 19922 33640 22066
rect 33888 21962 33916 22578
rect 33876 21956 33928 21962
rect 33876 21898 33928 21904
rect 33888 21865 33916 21898
rect 33874 21856 33930 21865
rect 33874 21791 33930 21800
rect 33980 21146 34008 26046
rect 34256 23254 34284 26302
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26200 37058 27000
rect 37646 26330 37702 27000
rect 37646 26302 37872 26330
rect 37646 26200 37702 26302
rect 34334 24712 34390 24721
rect 34334 24647 34390 24656
rect 34348 23662 34376 24647
rect 34440 23662 34468 26200
rect 34794 25936 34850 25945
rect 34794 25871 34850 25880
rect 34704 25424 34756 25430
rect 34704 25366 34756 25372
rect 34612 25356 34664 25362
rect 34612 25298 34664 25304
rect 34624 23730 34652 25298
rect 34612 23724 34664 23730
rect 34612 23666 34664 23672
rect 34336 23656 34388 23662
rect 34336 23598 34388 23604
rect 34428 23656 34480 23662
rect 34428 23598 34480 23604
rect 34244 23248 34296 23254
rect 34244 23190 34296 23196
rect 34336 23112 34388 23118
rect 34336 23054 34388 23060
rect 34348 22778 34376 23054
rect 34336 22772 34388 22778
rect 34336 22714 34388 22720
rect 34428 22704 34480 22710
rect 34428 22646 34480 22652
rect 34336 22568 34388 22574
rect 34336 22510 34388 22516
rect 34348 21622 34376 22510
rect 34440 22166 34468 22646
rect 34716 22642 34744 25366
rect 34808 23186 34836 25871
rect 35084 24562 35112 26200
rect 35256 26036 35308 26042
rect 35256 25978 35308 25984
rect 35084 24534 35204 24562
rect 35072 24404 35124 24410
rect 35072 24346 35124 24352
rect 34886 24304 34942 24313
rect 34886 24239 34942 24248
rect 34900 24206 34928 24239
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 34980 23316 35032 23322
rect 34980 23258 35032 23264
rect 34796 23180 34848 23186
rect 34796 23122 34848 23128
rect 34992 23050 35020 23258
rect 35084 23225 35112 24346
rect 35070 23216 35126 23225
rect 35070 23151 35126 23160
rect 35084 23118 35112 23151
rect 35072 23112 35124 23118
rect 35072 23054 35124 23060
rect 35176 23050 35204 24534
rect 34980 23044 35032 23050
rect 34980 22986 35032 22992
rect 35164 23044 35216 23050
rect 35164 22986 35216 22992
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 34428 22160 34480 22166
rect 34428 22102 34480 22108
rect 35268 22098 35296 25978
rect 35624 24948 35676 24954
rect 35624 24890 35676 24896
rect 35636 23594 35664 24890
rect 35728 24818 35756 26200
rect 36084 25968 36136 25974
rect 36084 25910 36136 25916
rect 35900 25560 35952 25566
rect 35900 25502 35952 25508
rect 35990 25528 36046 25537
rect 35806 25256 35862 25265
rect 35806 25191 35862 25200
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 35820 24206 35848 25191
rect 35808 24200 35860 24206
rect 35808 24142 35860 24148
rect 35808 24064 35860 24070
rect 35808 24006 35860 24012
rect 35716 23724 35768 23730
rect 35716 23666 35768 23672
rect 35624 23588 35676 23594
rect 35624 23530 35676 23536
rect 35728 23186 35756 23666
rect 35820 23662 35848 24006
rect 35912 23730 35940 25502
rect 35990 25463 36046 25472
rect 36004 24070 36032 25463
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 35808 23656 35860 23662
rect 35808 23598 35860 23604
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 35544 22953 35572 23054
rect 35900 22976 35952 22982
rect 35530 22944 35586 22953
rect 35900 22918 35952 22924
rect 35530 22879 35586 22888
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 34612 21956 34664 21962
rect 34612 21898 34664 21904
rect 34336 21616 34388 21622
rect 34334 21584 34336 21593
rect 34388 21584 34390 21593
rect 34334 21519 34390 21528
rect 34624 21350 34652 21898
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 34612 21344 34664 21350
rect 34612 21286 34664 21292
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 34336 20936 34388 20942
rect 34336 20878 34388 20884
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33600 19916 33652 19922
rect 33600 19858 33652 19864
rect 33138 19816 33194 19825
rect 33138 19751 33194 19760
rect 33152 19446 33180 19751
rect 33140 19440 33192 19446
rect 33140 19382 33192 19388
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32678 17504 32734 17513
rect 32678 17439 32734 17448
rect 32864 17060 32916 17066
rect 32864 17002 32916 17008
rect 32586 16008 32642 16017
rect 32586 15943 32642 15952
rect 32876 13841 32904 17002
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32862 13832 32918 13841
rect 32862 13767 32918 13776
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32220 13252 32272 13258
rect 32220 13194 32272 13200
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 31772 12406 31892 12434
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31404 9178 31432 11018
rect 31392 9172 31444 9178
rect 31392 9114 31444 9120
rect 29092 5296 29144 5302
rect 29144 5244 29224 5250
rect 29092 5238 29224 5244
rect 29104 5222 29224 5238
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 29104 2650 29132 5034
rect 29196 3670 29224 5222
rect 31772 5166 31800 12406
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 33336 6769 33364 19110
rect 33704 13977 33732 20402
rect 34348 20369 34376 20878
rect 34334 20360 34390 20369
rect 34334 20295 34390 20304
rect 33784 20256 33836 20262
rect 33784 20198 33836 20204
rect 33796 17785 33824 20198
rect 34348 20058 34376 20295
rect 34520 20256 34572 20262
rect 34520 20198 34572 20204
rect 34336 20052 34388 20058
rect 34336 19994 34388 20000
rect 33782 17776 33838 17785
rect 33782 17711 33838 17720
rect 34532 17066 34560 20198
rect 34520 17060 34572 17066
rect 34520 17002 34572 17008
rect 34716 14385 34744 21626
rect 35544 21622 35572 22879
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 35532 21616 35584 21622
rect 35532 21558 35584 21564
rect 34888 21548 34940 21554
rect 34888 21490 34940 21496
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 34900 19718 34928 21490
rect 35360 20913 35388 21490
rect 35346 20904 35402 20913
rect 35256 20868 35308 20874
rect 35530 20904 35586 20913
rect 35346 20839 35402 20848
rect 35440 20868 35492 20874
rect 35256 20810 35308 20816
rect 35530 20839 35586 20848
rect 35440 20810 35492 20816
rect 35072 20800 35124 20806
rect 35072 20742 35124 20748
rect 34980 20596 35032 20602
rect 34980 20538 35032 20544
rect 34992 20330 35020 20538
rect 34980 20324 35032 20330
rect 34980 20266 35032 20272
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34702 14376 34758 14385
rect 34702 14311 34758 14320
rect 33690 13968 33746 13977
rect 33690 13903 33746 13912
rect 34900 10470 34928 19654
rect 34888 10464 34940 10470
rect 34888 10406 34940 10412
rect 35084 10033 35112 20742
rect 35164 20324 35216 20330
rect 35164 20266 35216 20272
rect 35070 10024 35126 10033
rect 35070 9959 35126 9968
rect 35176 9489 35204 20266
rect 35268 20262 35296 20810
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 35256 20256 35308 20262
rect 35256 20198 35308 20204
rect 35268 18193 35296 20198
rect 35254 18184 35310 18193
rect 35254 18119 35310 18128
rect 35360 11898 35388 20266
rect 35452 20262 35480 20810
rect 35544 20602 35572 20839
rect 35532 20596 35584 20602
rect 35532 20538 35584 20544
rect 35636 20398 35664 22578
rect 35912 22438 35940 22918
rect 35992 22568 36044 22574
rect 35992 22510 36044 22516
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35716 21956 35768 21962
rect 35716 21898 35768 21904
rect 35900 21956 35952 21962
rect 35900 21898 35952 21904
rect 35624 20392 35676 20398
rect 35624 20334 35676 20340
rect 35728 20330 35756 21898
rect 35912 21457 35940 21898
rect 35898 21448 35954 21457
rect 35898 21383 35954 21392
rect 35716 20324 35768 20330
rect 35716 20266 35768 20272
rect 35440 20256 35492 20262
rect 35440 20198 35492 20204
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35162 9480 35218 9489
rect 35162 9415 35218 9424
rect 35452 9042 35480 20198
rect 36004 12345 36032 22510
rect 36096 22438 36124 25910
rect 36268 25628 36320 25634
rect 36268 25570 36320 25576
rect 36280 24290 36308 25570
rect 36188 24262 36308 24290
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 36188 21690 36216 24262
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 36280 22098 36308 22170
rect 36268 22092 36320 22098
rect 36268 22034 36320 22040
rect 36268 21888 36320 21894
rect 36268 21830 36320 21836
rect 36176 21684 36228 21690
rect 36176 21626 36228 21632
rect 36280 21554 36308 21830
rect 36372 21554 36400 26200
rect 37016 25786 37044 26200
rect 36544 25764 36596 25770
rect 37016 25758 37136 25786
rect 36544 25706 36596 25712
rect 36556 23866 36584 25706
rect 37002 25664 37058 25673
rect 37002 25599 37058 25608
rect 36636 24676 36688 24682
rect 36636 24618 36688 24624
rect 36544 23860 36596 23866
rect 36544 23802 36596 23808
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36464 23254 36492 23666
rect 36452 23248 36504 23254
rect 36452 23190 36504 23196
rect 36648 22710 36676 24618
rect 37016 24614 37044 25599
rect 36912 24608 36964 24614
rect 36912 24550 36964 24556
rect 37004 24608 37056 24614
rect 37004 24550 37056 24556
rect 36726 24168 36782 24177
rect 36726 24103 36782 24112
rect 36740 24070 36768 24103
rect 36728 24064 36780 24070
rect 36728 24006 36780 24012
rect 36924 23866 36952 24550
rect 36912 23860 36964 23866
rect 36912 23802 36964 23808
rect 36912 23724 36964 23730
rect 36912 23666 36964 23672
rect 36924 23254 36952 23666
rect 37108 23322 37136 25758
rect 37462 25392 37518 25401
rect 37462 25327 37518 25336
rect 37372 24132 37424 24138
rect 37372 24074 37424 24080
rect 37280 24064 37332 24070
rect 37280 24006 37332 24012
rect 37292 23338 37320 24006
rect 37004 23316 37056 23322
rect 37004 23258 37056 23264
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 37200 23310 37320 23338
rect 36912 23248 36964 23254
rect 36912 23190 36964 23196
rect 36728 23180 36780 23186
rect 36780 23140 36860 23168
rect 36728 23122 36780 23128
rect 36636 22704 36688 22710
rect 36636 22646 36688 22652
rect 36728 22636 36780 22642
rect 36728 22578 36780 22584
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36740 21418 36768 22578
rect 36832 21690 36860 23140
rect 37016 23118 37044 23258
rect 37004 23112 37056 23118
rect 37004 23054 37056 23060
rect 37200 22982 37228 23310
rect 37280 23248 37332 23254
rect 37280 23190 37332 23196
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37292 22545 37320 23190
rect 37384 23050 37412 24074
rect 37476 23866 37504 25327
rect 37740 24744 37792 24750
rect 37740 24686 37792 24692
rect 37464 23860 37516 23866
rect 37464 23802 37516 23808
rect 37752 23730 37780 24686
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37464 23112 37516 23118
rect 37464 23054 37516 23060
rect 37372 23044 37424 23050
rect 37372 22986 37424 22992
rect 37384 22710 37412 22986
rect 37372 22704 37424 22710
rect 37372 22646 37424 22652
rect 37278 22536 37334 22545
rect 37278 22471 37334 22480
rect 36912 22432 36964 22438
rect 36912 22374 36964 22380
rect 36820 21684 36872 21690
rect 36820 21626 36872 21632
rect 36728 21412 36780 21418
rect 36728 21354 36780 21360
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36452 20868 36504 20874
rect 36452 20810 36504 20816
rect 35990 12336 36046 12345
rect 35990 12271 36046 12280
rect 35440 9036 35492 9042
rect 35440 8978 35492 8984
rect 36464 8945 36492 20810
rect 36544 20800 36596 20806
rect 36544 20742 36596 20748
rect 36556 9625 36584 20742
rect 36648 19417 36676 20878
rect 36634 19408 36690 19417
rect 36634 19343 36690 19352
rect 36542 9616 36598 9625
rect 36542 9551 36598 9560
rect 36450 8936 36506 8945
rect 36450 8871 36506 8880
rect 36740 8401 36768 21354
rect 36924 21350 36952 22374
rect 37476 22094 37504 23054
rect 37556 23044 37608 23050
rect 37556 22986 37608 22992
rect 37384 22066 37504 22094
rect 37096 22024 37148 22030
rect 37016 21972 37096 21978
rect 37016 21966 37148 21972
rect 37016 21950 37136 21966
rect 36912 21344 36964 21350
rect 36912 21286 36964 21292
rect 36726 8392 36782 8401
rect 36726 8327 36782 8336
rect 37016 7449 37044 21950
rect 37096 21888 37148 21894
rect 37096 21830 37148 21836
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 37108 20806 37136 21830
rect 37096 20800 37148 20806
rect 37096 20742 37148 20748
rect 37108 13297 37136 20742
rect 37200 18426 37228 21830
rect 37384 21146 37412 22066
rect 37372 21140 37424 21146
rect 37372 21082 37424 21088
rect 37568 19514 37596 22986
rect 37648 22976 37700 22982
rect 37648 22918 37700 22924
rect 37556 19508 37608 19514
rect 37556 19450 37608 19456
rect 37188 18420 37240 18426
rect 37188 18362 37240 18368
rect 37660 13433 37688 22918
rect 37844 22658 37872 26302
rect 38290 26200 38346 27000
rect 38750 26208 38806 26217
rect 38304 24206 38332 26200
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 40866 26200 40922 27000
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26330 45430 27000
rect 45374 26302 45508 26330
rect 45374 26200 45430 26302
rect 38750 26143 38806 26152
rect 38474 25800 38530 25809
rect 38474 25735 38530 25744
rect 38384 24812 38436 24818
rect 38384 24754 38436 24760
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38304 23594 38332 24142
rect 38292 23588 38344 23594
rect 38292 23530 38344 23536
rect 38292 23044 38344 23050
rect 38292 22986 38344 22992
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37844 22630 37964 22658
rect 37832 22568 37884 22574
rect 37832 22510 37884 22516
rect 37740 22024 37792 22030
rect 37740 21966 37792 21972
rect 37752 21434 37780 21966
rect 37844 21690 37872 22510
rect 37936 22030 37964 22630
rect 38304 22234 38332 22986
rect 38396 22438 38424 24754
rect 38488 23118 38516 25735
rect 38660 25696 38712 25702
rect 38660 25638 38712 25644
rect 38672 24274 38700 25638
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 38764 23866 38792 26143
rect 38948 24206 38976 26200
rect 39118 25120 39174 25129
rect 39118 25055 39174 25064
rect 38936 24200 38988 24206
rect 38936 24142 38988 24148
rect 38752 23860 38804 23866
rect 38752 23802 38804 23808
rect 38476 23112 38528 23118
rect 38476 23054 38528 23060
rect 38936 23112 38988 23118
rect 38936 23054 38988 23060
rect 38384 22432 38436 22438
rect 38384 22374 38436 22380
rect 38292 22228 38344 22234
rect 38292 22170 38344 22176
rect 37924 22024 37976 22030
rect 37924 21966 37976 21972
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 38304 21622 38332 21966
rect 38292 21616 38344 21622
rect 38292 21558 38344 21564
rect 37752 21406 37872 21434
rect 37844 21350 37872 21406
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37844 18737 37872 21286
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38948 19281 38976 23054
rect 39132 22982 39160 25055
rect 39304 24608 39356 24614
rect 39304 24550 39356 24556
rect 39316 24410 39344 24550
rect 39304 24404 39356 24410
rect 39304 24346 39356 24352
rect 39212 24200 39264 24206
rect 39212 24142 39264 24148
rect 39224 23866 39252 24142
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 39120 22976 39172 22982
rect 39120 22918 39172 22924
rect 39224 22094 39252 23666
rect 39592 23662 39620 26200
rect 39764 25832 39816 25838
rect 39764 25774 39816 25780
rect 39580 23656 39632 23662
rect 39580 23598 39632 23604
rect 39776 23118 39804 25774
rect 39856 25084 39908 25090
rect 39856 25026 39908 25032
rect 39764 23112 39816 23118
rect 39764 23054 39816 23060
rect 39580 23044 39632 23050
rect 39580 22986 39632 22992
rect 39488 22704 39540 22710
rect 39488 22646 39540 22652
rect 39500 22234 39528 22646
rect 39488 22228 39540 22234
rect 39488 22170 39540 22176
rect 39224 22066 39344 22094
rect 38934 19272 38990 19281
rect 38934 19207 38990 19216
rect 37830 18728 37886 18737
rect 37830 18663 37886 18672
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37646 13424 37702 13433
rect 37646 13359 37702 13368
rect 37094 13288 37150 13297
rect 37094 13223 37150 13232
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 39316 11762 39344 22066
rect 39592 20534 39620 22986
rect 39776 22794 39804 23054
rect 39868 22982 39896 25026
rect 40040 25016 40092 25022
rect 40040 24958 40092 24964
rect 40052 24410 40080 24958
rect 40132 24880 40184 24886
rect 40132 24822 40184 24828
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 40144 23730 40172 24822
rect 40236 24188 40264 26200
rect 40408 25900 40460 25906
rect 40408 25842 40460 25848
rect 40316 24200 40368 24206
rect 40236 24160 40316 24188
rect 40316 24142 40368 24148
rect 40420 23730 40448 25842
rect 40776 24064 40828 24070
rect 40776 24006 40828 24012
rect 40788 23798 40816 24006
rect 40776 23792 40828 23798
rect 40776 23734 40828 23740
rect 39948 23724 40000 23730
rect 39948 23666 40000 23672
rect 40132 23724 40184 23730
rect 40132 23666 40184 23672
rect 40408 23724 40460 23730
rect 40408 23666 40460 23672
rect 39856 22976 39908 22982
rect 39856 22918 39908 22924
rect 39960 22794 39988 23666
rect 40144 23474 40172 23666
rect 40224 23520 40276 23526
rect 40144 23468 40224 23474
rect 40144 23462 40276 23468
rect 40144 23446 40264 23462
rect 40880 23254 40908 26200
rect 41524 24290 41552 26200
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 41524 24262 41644 24290
rect 41616 24206 41644 24262
rect 41236 24200 41288 24206
rect 41236 24142 41288 24148
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 41604 24200 41656 24206
rect 41604 24142 41656 24148
rect 42616 24200 42668 24206
rect 42616 24142 42668 24148
rect 41248 23798 41276 24142
rect 41236 23792 41288 23798
rect 41236 23734 41288 23740
rect 40960 23656 41012 23662
rect 40960 23598 41012 23604
rect 41052 23656 41104 23662
rect 41052 23598 41104 23604
rect 40868 23248 40920 23254
rect 40868 23190 40920 23196
rect 40868 23112 40920 23118
rect 40868 23054 40920 23060
rect 39776 22766 39896 22794
rect 39960 22778 40080 22794
rect 39960 22772 40092 22778
rect 39960 22766 40040 22772
rect 39764 22432 39816 22438
rect 39764 22374 39816 22380
rect 39580 20528 39632 20534
rect 39580 20470 39632 20476
rect 39776 19310 39804 22374
rect 39868 22098 39896 22766
rect 40040 22714 40092 22720
rect 40880 22506 40908 23054
rect 40868 22500 40920 22506
rect 40868 22442 40920 22448
rect 39856 22092 39908 22098
rect 39856 22034 39908 22040
rect 40972 20466 41000 23598
rect 41064 23526 41092 23598
rect 41052 23520 41104 23526
rect 41052 23462 41104 23468
rect 41144 23112 41196 23118
rect 41144 23054 41196 23060
rect 41156 22778 41184 23054
rect 41144 22772 41196 22778
rect 41144 22714 41196 22720
rect 40960 20460 41012 20466
rect 40960 20402 41012 20408
rect 39764 19304 39816 19310
rect 39764 19246 39816 19252
rect 41524 12889 41552 24142
rect 42432 24132 42484 24138
rect 42432 24074 42484 24080
rect 42524 24132 42576 24138
rect 42524 24074 42576 24080
rect 42444 23866 42472 24074
rect 42432 23860 42484 23866
rect 42432 23802 42484 23808
rect 41972 22976 42024 22982
rect 41972 22918 42024 22924
rect 41984 19786 42012 22918
rect 41972 19780 42024 19786
rect 41972 19722 42024 19728
rect 42536 18698 42564 24074
rect 42628 23866 42656 24142
rect 43456 23866 43484 26200
rect 43536 24336 43588 24342
rect 43536 24278 43588 24284
rect 42616 23860 42668 23866
rect 42616 23802 42668 23808
rect 43444 23860 43496 23866
rect 43444 23802 43496 23808
rect 43444 23588 43496 23594
rect 43444 23530 43496 23536
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42524 18692 42576 18698
rect 42524 18634 42576 18640
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 43456 14958 43484 23530
rect 43548 16182 43576 24278
rect 43904 24064 43956 24070
rect 43904 24006 43956 24012
rect 43720 23520 43772 23526
rect 43720 23462 43772 23468
rect 43732 18630 43760 23462
rect 43916 22710 43944 24006
rect 44100 23712 44128 26200
rect 44744 24410 44772 26200
rect 44732 24404 44784 24410
rect 44732 24346 44784 24352
rect 44744 24206 44772 24346
rect 45480 24290 45508 26302
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26330 48650 27000
rect 48594 26302 48912 26330
rect 48594 26200 48650 26302
rect 45834 24848 45890 24857
rect 45834 24783 45890 24792
rect 45480 24262 45600 24290
rect 45572 24206 45600 24262
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 45284 24064 45336 24070
rect 45284 24006 45336 24012
rect 44180 23724 44232 23730
rect 44100 23684 44180 23712
rect 44180 23666 44232 23672
rect 43904 22704 43956 22710
rect 43904 22646 43956 22652
rect 43720 18624 43772 18630
rect 43720 18566 43772 18572
rect 43536 16176 43588 16182
rect 43536 16118 43588 16124
rect 45296 15910 45324 24006
rect 45572 23866 45600 24142
rect 45560 23860 45612 23866
rect 45560 23802 45612 23808
rect 45466 23080 45522 23089
rect 45466 23015 45522 23024
rect 45480 17610 45508 23015
rect 45848 19242 45876 24783
rect 46032 24206 46060 26200
rect 46020 24200 46072 24206
rect 46020 24142 46072 24148
rect 46202 23760 46258 23769
rect 46676 23730 46704 26200
rect 47320 24206 47348 26200
rect 47964 24206 47992 26200
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 47952 24200 48004 24206
rect 47952 24142 48004 24148
rect 47032 24064 47084 24070
rect 47032 24006 47084 24012
rect 46202 23695 46258 23704
rect 46664 23724 46716 23730
rect 45836 19236 45888 19242
rect 45836 19178 45888 19184
rect 45468 17604 45520 17610
rect 45468 17546 45520 17552
rect 45284 15904 45336 15910
rect 45284 15846 45336 15852
rect 43444 14952 43496 14958
rect 43444 14894 43496 14900
rect 46216 14890 46244 23695
rect 46664 23666 46716 23672
rect 46940 23520 46992 23526
rect 46940 23462 46992 23468
rect 46846 21992 46902 22001
rect 46846 21927 46902 21936
rect 46860 20942 46888 21927
rect 46848 20936 46900 20942
rect 46848 20878 46900 20884
rect 46952 15978 46980 23462
rect 47044 17542 47072 24006
rect 47320 23866 47348 24142
rect 48596 24064 48648 24070
rect 48596 24006 48648 24012
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47584 21548 47636 21554
rect 47584 21490 47636 21496
rect 47596 21350 47624 21490
rect 47584 21344 47636 21350
rect 47584 21286 47636 21292
rect 47032 17536 47084 17542
rect 47032 17478 47084 17484
rect 46940 15972 46992 15978
rect 46940 15914 46992 15920
rect 46204 14884 46256 14890
rect 46204 14826 46256 14832
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 41510 12880 41566 12889
rect 41510 12815 41566 12824
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 39304 11756 39356 11762
rect 39304 11698 39356 11704
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 47596 11150 47624 21286
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 48608 14822 48636 24006
rect 48884 23730 48912 26302
rect 48872 23724 48924 23730
rect 48872 23666 48924 23672
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48700 22574 48728 23462
rect 48688 22568 48740 22574
rect 48688 22510 48740 22516
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 48596 14816 48648 14822
rect 48596 14758 48648 14764
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47584 11144 47636 11150
rect 47584 11086 47636 11092
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 37002 7440 37058 7449
rect 37002 7375 37058 7384
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 33322 6760 33378 6769
rect 33322 6695 33378 6704
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 31760 5160 31812 5166
rect 31760 5102 31812 5108
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 29656 4758 29684 5102
rect 29644 4752 29696 4758
rect 29644 4694 29696 4700
rect 32508 3738 32536 5102
rect 32864 5092 32916 5098
rect 32864 5034 32916 5040
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 29184 3664 29236 3670
rect 29184 3606 29236 3612
rect 32876 2650 32904 5034
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 41420 3732 41472 3738
rect 41420 3674 41472 3680
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 25424 800 25452 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 3402
rect 41432 800 41460 3674
rect 44088 3664 44140 3670
rect 44088 3606 44140 3612
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 44100 800 44128 3606
rect 46756 3596 46808 3602
rect 46756 3538 46808 3544
rect 46768 800 46796 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 3470
rect 28184 734 28396 762
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 1582 24284 1584 24304
rect 1584 24284 1636 24304
rect 1636 24284 1638 24304
rect 1582 24248 1638 24284
rect 1766 24148 1768 24168
rect 1768 24148 1820 24168
rect 1820 24148 1822 24168
rect 1766 24112 1822 24148
rect 1306 20712 1362 20768
rect 1858 20440 1914 20496
rect 1674 19624 1730 19680
rect 1398 17856 1454 17912
rect 1214 17040 1270 17096
rect 1122 16360 1178 16416
rect 1122 16088 1178 16144
rect 1122 15000 1178 15056
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 938 10668 994 10704
rect 938 10648 940 10668
rect 940 10648 992 10668
rect 992 10648 994 10668
rect 1122 13368 1178 13424
rect 1766 13368 1822 13424
rect 1582 11092 1584 11112
rect 1584 11092 1636 11112
rect 1636 11092 1638 11112
rect 1582 11056 1638 11092
rect 1766 12144 1822 12200
rect 2042 17448 2098 17504
rect 2042 13776 2098 13832
rect 1490 9596 1492 9616
rect 1492 9596 1544 9616
rect 1544 9596 1546 9616
rect 1490 9560 1546 9596
rect 1858 11600 1914 11656
rect 1858 10920 1914 10976
rect 1858 10668 1914 10704
rect 1858 10648 1860 10668
rect 1860 10648 1912 10668
rect 1912 10648 1914 10668
rect 2042 11056 2098 11112
rect 3146 25200 3202 25256
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2778 24384 2834 24440
rect 3882 25608 3938 25664
rect 3698 24792 3754 24848
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2686 21528 2742 21584
rect 1306 6024 1362 6080
rect 1582 5616 1638 5672
rect 1306 5208 1362 5264
rect 1582 4800 1638 4856
rect 2778 21120 2834 21176
rect 3514 22480 3570 22536
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3422 21528 3478 21584
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 3330 19896 3386 19952
rect 2686 19080 2742 19136
rect 2594 18808 2650 18864
rect 2502 12280 2558 12336
rect 2410 11892 2466 11928
rect 2410 11872 2412 11892
rect 2412 11872 2464 11892
rect 2464 11872 2466 11892
rect 2410 10376 2466 10432
rect 2318 8064 2374 8120
rect 2962 19488 3018 19544
rect 3330 19236 3386 19272
rect 3330 19216 3332 19236
rect 3332 19216 3384 19236
rect 3384 19216 3386 19236
rect 3974 24656 4030 24712
rect 4066 23976 4122 24032
rect 3974 23568 4030 23624
rect 4250 24792 4306 24848
rect 3882 23160 3938 23216
rect 4066 23024 4122 23080
rect 4066 22752 4122 22808
rect 3974 22616 4030 22672
rect 3698 21936 3754 21992
rect 3790 21664 3846 21720
rect 3606 20848 3662 20904
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18672 2926 18728
rect 2778 18264 2834 18320
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 3330 17720 3386 17776
rect 3606 20168 3662 20224
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 3606 19372 3662 19408
rect 3606 19352 3608 19372
rect 3608 19352 3660 19372
rect 3660 19352 3662 19372
rect 3606 19080 3662 19136
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 3422 16632 3478 16688
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 3422 15408 3478 15464
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3238 12960 3294 13016
rect 3606 14476 3662 14512
rect 3606 14456 3608 14476
rect 3608 14456 3660 14476
rect 3660 14456 3662 14476
rect 3514 13912 3570 13968
rect 3330 12552 3386 12608
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 3238 12180 3240 12200
rect 3240 12180 3292 12200
rect 3292 12180 3294 12200
rect 3238 12144 3294 12180
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2870 10784 2926 10840
rect 2778 9288 2834 9344
rect 2778 7792 2834 7848
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2962 9988 3018 10024
rect 2962 9968 2964 9988
rect 2964 9968 3016 9988
rect 3016 9968 3018 9988
rect 3606 13504 3662 13560
rect 3606 12552 3662 12608
rect 3606 11328 3662 11384
rect 3698 11192 3754 11248
rect 3422 10512 3478 10568
rect 3330 9596 3332 9616
rect 3332 9596 3384 9616
rect 3384 9596 3386 9616
rect 3330 9560 3386 9596
rect 3606 10104 3662 10160
rect 3514 9696 3570 9752
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3146 8880 3202 8936
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3238 7384 3294 7440
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3146 6704 3202 6760
rect 2870 6568 2926 6624
rect 3146 6296 3202 6352
rect 2870 6160 2926 6216
rect 1214 3984 1270 4040
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3422 9444 3478 9480
rect 3422 9424 3424 9444
rect 3424 9424 3476 9444
rect 3476 9424 3478 9444
rect 3790 10804 3846 10840
rect 3790 10784 3792 10804
rect 3792 10784 3844 10804
rect 3844 10784 3846 10804
rect 4158 18944 4214 19000
rect 4066 17620 4068 17640
rect 4068 17620 4120 17640
rect 4120 17620 4122 17640
rect 4066 17584 4122 17620
rect 4158 15952 4214 16008
rect 4066 12844 4122 12880
rect 4066 12824 4068 12844
rect 4068 12824 4120 12844
rect 4120 12824 4122 12844
rect 4066 12436 4122 12472
rect 4066 12416 4068 12436
rect 4068 12416 4120 12436
rect 4120 12416 4122 12436
rect 4066 12280 4122 12336
rect 3974 9560 4030 9616
rect 3882 9152 3938 9208
rect 3882 9016 3938 9072
rect 4618 22344 4674 22400
rect 4434 15544 4490 15600
rect 4342 15308 4344 15328
rect 4344 15308 4396 15328
rect 4396 15308 4398 15328
rect 4342 15272 4398 15308
rect 4434 13912 4490 13968
rect 4434 13232 4490 13288
rect 4342 12280 4398 12336
rect 4434 12008 4490 12064
rect 5170 21392 5226 21448
rect 4710 15816 4766 15872
rect 4618 12688 4674 12744
rect 4526 9832 4582 9888
rect 4250 9460 4252 9480
rect 4252 9460 4304 9480
rect 4304 9460 4306 9480
rect 4250 9424 4306 9460
rect 4250 8900 4306 8936
rect 4250 8880 4252 8900
rect 4252 8880 4304 8900
rect 4304 8880 4306 8900
rect 4342 7656 4398 7712
rect 4250 6432 4306 6488
rect 3974 6296 4030 6352
rect 4158 6316 4214 6352
rect 4158 6296 4160 6316
rect 4160 6296 4212 6316
rect 4212 6296 4214 6316
rect 4158 6060 4160 6080
rect 4160 6060 4212 6080
rect 4212 6060 4214 6080
rect 4158 6024 4214 6060
rect 4158 5752 4214 5808
rect 3330 4664 3386 4720
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 3596 1362 3632
rect 5998 21936 6054 21992
rect 5630 21800 5686 21856
rect 5906 21256 5962 21312
rect 5814 21140 5870 21176
rect 5814 21120 5816 21140
rect 5816 21120 5868 21140
rect 5868 21120 5870 21140
rect 5906 20576 5962 20632
rect 5446 18536 5502 18592
rect 5354 18128 5410 18184
rect 5170 17856 5226 17912
rect 4710 10104 4766 10160
rect 5170 15680 5226 15736
rect 4894 13640 4950 13696
rect 4986 13096 5042 13152
rect 4894 12008 4950 12064
rect 4802 8472 4858 8528
rect 4710 7928 4766 7984
rect 4618 7520 4674 7576
rect 4526 7248 4582 7304
rect 4894 8200 4950 8256
rect 5630 17040 5686 17096
rect 5446 16496 5502 16552
rect 5630 16244 5686 16280
rect 5630 16224 5632 16244
rect 5632 16224 5684 16244
rect 5684 16224 5686 16244
rect 5906 18808 5962 18864
rect 5814 15816 5870 15872
rect 5262 13640 5318 13696
rect 5538 13776 5594 13832
rect 5354 12824 5410 12880
rect 5630 12280 5686 12336
rect 5354 12008 5410 12064
rect 5538 10920 5594 10976
rect 5170 9016 5226 9072
rect 5998 17856 6054 17912
rect 6458 24928 6514 24984
rect 6458 22480 6514 22536
rect 7378 25472 7434 25528
rect 6826 23196 6828 23216
rect 6828 23196 6880 23216
rect 6880 23196 6882 23216
rect 6826 23160 6882 23196
rect 6918 22636 6974 22672
rect 6918 22616 6920 22636
rect 6920 22616 6972 22636
rect 6972 22616 6974 22636
rect 6274 19508 6330 19544
rect 6274 19488 6276 19508
rect 6276 19488 6328 19508
rect 6328 19488 6330 19508
rect 6090 16224 6146 16280
rect 5998 15544 6054 15600
rect 5998 15020 6054 15056
rect 5998 15000 6000 15020
rect 6000 15000 6052 15020
rect 6052 15000 6054 15020
rect 6366 16768 6422 16824
rect 6090 12860 6092 12880
rect 6092 12860 6144 12880
rect 6144 12860 6146 12880
rect 6090 12824 6146 12860
rect 7378 22344 7434 22400
rect 6918 20304 6974 20360
rect 6550 19352 6606 19408
rect 7010 18400 7066 18456
rect 6366 15564 6422 15600
rect 6366 15544 6368 15564
rect 6368 15544 6420 15564
rect 6420 15544 6422 15564
rect 6274 12824 6330 12880
rect 6366 12300 6422 12336
rect 6366 12280 6368 12300
rect 6368 12280 6420 12300
rect 6420 12280 6422 12300
rect 6550 12008 6606 12064
rect 7010 17620 7012 17640
rect 7012 17620 7064 17640
rect 7064 17620 7066 17640
rect 7010 17584 7066 17620
rect 7378 19760 7434 19816
rect 7286 18572 7288 18592
rect 7288 18572 7340 18592
rect 7340 18572 7342 18592
rect 7286 18536 7342 18572
rect 7102 16088 7158 16144
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 8114 23568 8170 23624
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7930 21392 7986 21448
rect 8114 20984 8170 21040
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8390 19896 8446 19952
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8298 19352 8354 19408
rect 8298 18708 8300 18728
rect 8300 18708 8352 18728
rect 8352 18708 8354 18728
rect 8298 18672 8354 18708
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7838 17992 7894 18048
rect 7930 17856 7986 17912
rect 8206 18264 8262 18320
rect 8114 18128 8170 18184
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7930 16940 7932 16960
rect 7932 16940 7984 16960
rect 7984 16940 7986 16960
rect 7930 16904 7986 16940
rect 8114 16652 8170 16688
rect 8114 16632 8116 16652
rect 8116 16632 8168 16652
rect 8168 16632 8170 16652
rect 7746 16360 7802 16416
rect 7562 15544 7618 15600
rect 7194 13096 7250 13152
rect 5814 9696 5870 9752
rect 5998 9696 6054 9752
rect 5906 9016 5962 9072
rect 6274 9696 6330 9752
rect 6274 7112 6330 7168
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 6734 8200 6790 8256
rect 7010 9596 7012 9616
rect 7012 9596 7064 9616
rect 7064 9596 7066 9616
rect 7010 9560 7066 9596
rect 6918 9324 6920 9344
rect 6920 9324 6972 9344
rect 6972 9324 6974 9344
rect 6918 9288 6974 9324
rect 8206 14320 8262 14376
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7378 12008 7434 12064
rect 7286 11192 7342 11248
rect 7378 10376 7434 10432
rect 6826 7284 6828 7304
rect 6828 7284 6880 7304
rect 6880 7284 6882 7304
rect 6826 7248 6882 7284
rect 6918 6840 6974 6896
rect 9586 25200 9642 25256
rect 9310 23432 9366 23488
rect 9310 22072 9366 22128
rect 8574 18128 8630 18184
rect 8850 19352 8906 19408
rect 8850 16768 8906 16824
rect 8482 15816 8538 15872
rect 8482 14612 8538 14648
rect 8482 14592 8484 14612
rect 8484 14592 8536 14612
rect 8536 14592 8538 14612
rect 9494 22208 9550 22264
rect 9402 19896 9458 19952
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 8114 11328 8170 11384
rect 7378 7404 7434 7440
rect 7378 7384 7380 7404
rect 7380 7384 7432 7404
rect 7432 7384 7434 7404
rect 7194 6996 7250 7032
rect 7194 6976 7196 6996
rect 7196 6976 7248 6996
rect 7248 6976 7250 6996
rect 7010 6568 7066 6624
rect 6918 6432 6974 6488
rect 3698 4392 3754 4448
rect 1306 3576 1308 3596
rect 1308 3576 1360 3596
rect 1360 3576 1362 3596
rect 1306 2760 1362 2816
rect 1306 2352 1362 2408
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 4066 3168 4122 3224
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 8850 14320 8906 14376
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8298 8472 8354 8528
rect 8114 8372 8116 8392
rect 8116 8372 8168 8392
rect 8168 8372 8170 8392
rect 8114 8336 8170 8372
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7838 5616 7894 5672
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 8298 4664 8354 4720
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 8482 8200 8538 8256
rect 8666 7520 8722 7576
rect 8482 6432 8538 6488
rect 10046 23704 10102 23760
rect 9770 22888 9826 22944
rect 9954 20576 10010 20632
rect 9586 18808 9642 18864
rect 9678 18672 9734 18728
rect 9402 16768 9458 16824
rect 9402 15952 9458 16008
rect 9770 18536 9826 18592
rect 9586 17992 9642 18048
rect 9678 17856 9734 17912
rect 9586 15816 9642 15872
rect 9954 16360 10010 16416
rect 8942 9696 8998 9752
rect 9586 13812 9588 13832
rect 9588 13812 9640 13832
rect 9640 13812 9642 13832
rect 9586 13776 9642 13812
rect 9310 8472 9366 8528
rect 9402 7948 9458 7984
rect 9402 7928 9404 7948
rect 9404 7928 9456 7948
rect 9456 7928 9458 7948
rect 9770 14592 9826 14648
rect 9770 11464 9826 11520
rect 9770 10956 9772 10976
rect 9772 10956 9824 10976
rect 9824 10956 9826 10976
rect 9770 10920 9826 10956
rect 10138 19216 10194 19272
rect 11150 23840 11206 23896
rect 11058 22772 11114 22808
rect 11058 22752 11060 22772
rect 11060 22752 11112 22772
rect 11112 22752 11114 22772
rect 10690 21936 10746 21992
rect 10506 21664 10562 21720
rect 10506 21256 10562 21312
rect 10414 20984 10470 21040
rect 11058 22208 11114 22264
rect 11058 21664 11114 21720
rect 10966 21428 10968 21448
rect 10968 21428 11020 21448
rect 11020 21428 11022 21448
rect 10598 20712 10654 20768
rect 10506 20576 10562 20632
rect 10966 21392 11022 21428
rect 11794 22752 11850 22808
rect 11702 21800 11758 21856
rect 11150 21256 11206 21312
rect 10690 19624 10746 19680
rect 10322 18128 10378 18184
rect 10230 17312 10286 17368
rect 11150 19352 11206 19408
rect 10690 19080 10746 19136
rect 10598 18672 10654 18728
rect 10874 19080 10930 19136
rect 10690 18264 10746 18320
rect 10598 17992 10654 18048
rect 10874 17856 10930 17912
rect 10138 15136 10194 15192
rect 10138 14320 10194 14376
rect 10046 13640 10102 13696
rect 10598 16768 10654 16824
rect 10506 15952 10562 16008
rect 10690 14728 10746 14784
rect 9862 9696 9918 9752
rect 9678 9016 9734 9072
rect 9678 6976 9734 7032
rect 9862 8200 9918 8256
rect 9862 8064 9918 8120
rect 9862 7384 9918 7440
rect 10230 12960 10286 13016
rect 10046 8064 10102 8120
rect 12070 24384 12126 24440
rect 11978 24248 12034 24304
rect 11518 19896 11574 19952
rect 11518 19488 11574 19544
rect 11150 18264 11206 18320
rect 11150 17992 11206 18048
rect 11058 17448 11114 17504
rect 11058 16224 11114 16280
rect 10966 15816 11022 15872
rect 10966 14728 11022 14784
rect 10506 11736 10562 11792
rect 10506 11192 10562 11248
rect 10966 13796 11022 13832
rect 10966 13776 10968 13796
rect 10968 13776 11020 13796
rect 11020 13776 11022 13796
rect 10322 9560 10378 9616
rect 10322 8744 10378 8800
rect 10598 10648 10654 10704
rect 10506 9832 10562 9888
rect 10690 9696 10746 9752
rect 10690 9016 10746 9072
rect 10506 6724 10562 6760
rect 10506 6704 10508 6724
rect 10508 6704 10560 6724
rect 10560 6704 10562 6724
rect 11150 10784 11206 10840
rect 10966 9016 11022 9072
rect 11058 8628 11114 8664
rect 11058 8608 11060 8628
rect 11060 8608 11112 8628
rect 11112 8608 11114 8628
rect 11150 8472 11206 8528
rect 11610 18844 11612 18864
rect 11612 18844 11664 18864
rect 11664 18844 11666 18864
rect 11610 18808 11666 18844
rect 11610 18400 11666 18456
rect 11518 18264 11574 18320
rect 11426 16224 11482 16280
rect 11794 19080 11850 19136
rect 11794 18400 11850 18456
rect 11794 18300 11796 18320
rect 11796 18300 11848 18320
rect 11848 18300 11850 18320
rect 11794 18264 11850 18300
rect 11794 16940 11796 16960
rect 11796 16940 11848 16960
rect 11848 16940 11850 16960
rect 11794 16904 11850 16940
rect 11794 16360 11850 16416
rect 11426 14048 11482 14104
rect 11702 14456 11758 14512
rect 11610 13912 11666 13968
rect 11978 20440 12034 20496
rect 11978 19896 12034 19952
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12622 23024 12678 23080
rect 13174 22752 13230 22808
rect 13174 22480 13230 22536
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13634 26016 13690 26072
rect 12346 21528 12402 21584
rect 12530 21564 12532 21584
rect 12532 21564 12584 21584
rect 12584 21564 12586 21584
rect 12530 21528 12586 21564
rect 12346 20884 12348 20904
rect 12348 20884 12400 20904
rect 12400 20884 12402 20904
rect 12346 20848 12402 20884
rect 12530 20440 12586 20496
rect 12530 19896 12586 19952
rect 12346 19780 12402 19816
rect 12346 19760 12348 19780
rect 12348 19760 12400 19780
rect 12400 19760 12402 19780
rect 12162 19216 12218 19272
rect 12070 18400 12126 18456
rect 13358 21800 13414 21856
rect 13082 21664 13138 21720
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12806 21120 12862 21176
rect 13450 21120 13506 21176
rect 13726 24656 13782 24712
rect 13726 24112 13782 24168
rect 14830 24792 14886 24848
rect 14554 24520 14610 24576
rect 13818 22072 13874 22128
rect 13358 20340 13360 20360
rect 13360 20340 13412 20360
rect 13412 20340 13414 20360
rect 13358 20304 13414 20340
rect 12346 18944 12402 19000
rect 12346 17992 12402 18048
rect 11978 15136 12034 15192
rect 11978 14492 11980 14512
rect 11980 14492 12032 14512
rect 12032 14492 12034 14512
rect 11978 14456 12034 14492
rect 11978 12824 12034 12880
rect 11794 12552 11850 12608
rect 11794 12144 11850 12200
rect 12438 17448 12494 17504
rect 12346 16224 12402 16280
rect 12438 15680 12494 15736
rect 12162 15408 12218 15464
rect 12530 15544 12586 15600
rect 12254 14456 12310 14512
rect 12162 13932 12218 13968
rect 12162 13912 12164 13932
rect 12164 13912 12216 13932
rect 12216 13912 12218 13932
rect 11426 9288 11482 9344
rect 11334 8628 11390 8664
rect 11334 8608 11336 8628
rect 11336 8608 11388 8628
rect 11388 8608 11390 8628
rect 11334 7384 11390 7440
rect 10874 6568 10930 6624
rect 11978 11872 12034 11928
rect 11702 11736 11758 11792
rect 11610 8628 11666 8664
rect 11610 8608 11612 8628
rect 11612 8608 11664 8628
rect 11664 8608 11666 8628
rect 12070 11464 12126 11520
rect 12162 9832 12218 9888
rect 12346 8084 12402 8120
rect 12346 8064 12348 8084
rect 12348 8064 12400 8084
rect 12400 8064 12402 8084
rect 12806 20168 12862 20224
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12990 19760 13046 19816
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13358 18400 13414 18456
rect 12990 18164 12992 18184
rect 12992 18164 13044 18184
rect 13044 18164 13046 18184
rect 12990 18128 13046 18164
rect 14186 21392 14242 21448
rect 14186 20984 14242 21040
rect 13818 19488 13874 19544
rect 12806 17992 12862 18048
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12806 14592 12862 14648
rect 13910 18944 13966 19000
rect 13818 18400 13874 18456
rect 14094 18536 14150 18592
rect 13726 17176 13782 17232
rect 13818 16496 13874 16552
rect 13634 16360 13690 16416
rect 13818 16224 13874 16280
rect 13542 15308 13544 15328
rect 13544 15308 13596 15328
rect 13596 15308 13598 15328
rect 13542 15272 13598 15308
rect 12714 14320 12770 14376
rect 13358 14068 13414 14104
rect 13358 14048 13360 14068
rect 13360 14048 13412 14068
rect 13412 14048 13414 14068
rect 12898 13812 12900 13832
rect 12900 13812 12952 13832
rect 12952 13812 12954 13832
rect 12898 13776 12954 13812
rect 12806 13640 12862 13696
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13358 13504 13414 13560
rect 13910 15136 13966 15192
rect 13910 14884 13966 14920
rect 13910 14864 13912 14884
rect 13912 14864 13964 14884
rect 13964 14864 13966 14884
rect 13910 14184 13966 14240
rect 12714 12980 12770 13016
rect 12714 12960 12716 12980
rect 12716 12960 12768 12980
rect 12768 12960 12770 12980
rect 12990 12824 13046 12880
rect 13358 12960 13414 13016
rect 13542 12960 13598 13016
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12714 11328 12770 11384
rect 12530 8200 12586 8256
rect 12346 6976 12402 7032
rect 13174 11600 13230 11656
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13542 11328 13598 11384
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13266 9868 13268 9888
rect 13268 9868 13320 9888
rect 13320 9868 13322 9888
rect 13266 9832 13322 9868
rect 13266 9580 13322 9616
rect 13266 9560 13268 9580
rect 13268 9560 13320 9580
rect 13320 9560 13322 9580
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 14094 16632 14150 16688
rect 14094 15988 14096 16008
rect 14096 15988 14148 16008
rect 14148 15988 14150 16008
rect 14094 15952 14150 15988
rect 14094 15136 14150 15192
rect 14094 13096 14150 13152
rect 14186 12552 14242 12608
rect 14002 12008 14058 12064
rect 13174 9036 13230 9072
rect 13174 9016 13176 9036
rect 13176 9016 13228 9036
rect 13228 9016 13230 9036
rect 12806 8628 12862 8664
rect 12806 8608 12808 8628
rect 12808 8608 12860 8628
rect 12860 8608 12862 8628
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 13634 10920 13690 10976
rect 13358 7148 13360 7168
rect 13360 7148 13412 7168
rect 13412 7148 13414 7168
rect 13358 7112 13414 7148
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 13910 10784 13966 10840
rect 13910 8200 13966 8256
rect 13542 6160 13598 6216
rect 14186 11348 14242 11384
rect 14186 11328 14188 11348
rect 14188 11328 14240 11348
rect 14240 11328 14242 11348
rect 14554 24112 14610 24168
rect 14462 23160 14518 23216
rect 14830 23704 14886 23760
rect 14462 17720 14518 17776
rect 14462 16360 14518 16416
rect 15566 26152 15622 26208
rect 15290 23432 15346 23488
rect 16026 24384 16082 24440
rect 15658 23432 15714 23488
rect 14738 20848 14794 20904
rect 14830 18808 14886 18864
rect 14646 17584 14702 17640
rect 15106 20576 15162 20632
rect 16762 25880 16818 25936
rect 16578 25608 16634 25664
rect 16026 20304 16082 20360
rect 15474 18808 15530 18864
rect 14830 15680 14886 15736
rect 15014 15272 15070 15328
rect 15750 19896 15806 19952
rect 15658 19080 15714 19136
rect 15934 18536 15990 18592
rect 15750 17312 15806 17368
rect 15198 14320 15254 14376
rect 14554 12552 14610 12608
rect 14830 12552 14886 12608
rect 14646 12280 14702 12336
rect 14186 9560 14242 9616
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 15658 14048 15714 14104
rect 15382 12008 15438 12064
rect 15474 8608 15530 8664
rect 16026 16904 16082 16960
rect 16302 18028 16304 18048
rect 16304 18028 16356 18048
rect 16356 18028 16358 18048
rect 16302 17992 16358 18028
rect 16486 20032 16542 20088
rect 16762 25472 16818 25528
rect 16854 22888 16910 22944
rect 16394 17720 16450 17776
rect 16946 21428 16948 21448
rect 16948 21428 17000 21448
rect 17000 21428 17002 21448
rect 16946 21392 17002 21428
rect 17222 24792 17278 24848
rect 17958 26288 18014 26344
rect 17406 22752 17462 22808
rect 19246 26424 19302 26480
rect 17958 25880 18014 25936
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17958 23180 18014 23216
rect 17958 23160 17960 23180
rect 17960 23160 18012 23180
rect 18012 23160 18014 23180
rect 18878 24384 18934 24440
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 20074 24928 20130 24984
rect 19154 22888 19210 22944
rect 17130 21664 17186 21720
rect 18418 21800 18474 21856
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17038 19352 17094 19408
rect 17590 21256 17646 21312
rect 17866 21256 17922 21312
rect 18878 21936 18934 21992
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17682 20168 17738 20224
rect 17406 19216 17462 19272
rect 17314 18944 17370 19000
rect 16946 18572 16948 18592
rect 16948 18572 17000 18592
rect 17000 18572 17002 18592
rect 16946 18536 17002 18572
rect 16854 18148 16910 18184
rect 16854 18128 16856 18148
rect 16856 18128 16908 18148
rect 16908 18128 16910 18148
rect 15934 10532 15990 10568
rect 15934 10512 15936 10532
rect 15936 10512 15988 10532
rect 15988 10512 15990 10532
rect 16302 12008 16358 12064
rect 16762 16904 16818 16960
rect 17406 18400 17462 18456
rect 17314 16496 17370 16552
rect 17958 19916 18014 19952
rect 17958 19896 17960 19916
rect 17960 19896 18012 19916
rect 18012 19896 18014 19916
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18234 19372 18290 19408
rect 18234 19352 18236 19372
rect 18236 19352 18288 19372
rect 18288 19352 18290 19372
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18234 17584 18290 17640
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17222 15816 17278 15872
rect 16854 14456 16910 14512
rect 17222 14068 17278 14104
rect 17222 14048 17224 14068
rect 17224 14048 17276 14068
rect 17276 14048 17278 14068
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18050 13504 18106 13560
rect 18786 20576 18842 20632
rect 18694 20204 18696 20224
rect 18696 20204 18748 20224
rect 18748 20204 18750 20224
rect 18694 20168 18750 20204
rect 18418 17992 18474 18048
rect 18694 16768 18750 16824
rect 18418 13504 18474 13560
rect 16946 11600 17002 11656
rect 17498 11872 17554 11928
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 19798 23468 19800 23488
rect 19800 23468 19852 23488
rect 19852 23468 19854 23488
rect 19798 23432 19854 23468
rect 19982 22652 19984 22672
rect 19984 22652 20036 22672
rect 20036 22652 20038 22672
rect 19982 22616 20038 22652
rect 19614 22208 19670 22264
rect 21822 23976 21878 24032
rect 19522 21664 19578 21720
rect 19430 20748 19432 20768
rect 19432 20748 19484 20768
rect 19484 20748 19486 20768
rect 19430 20712 19486 20748
rect 19706 20324 19762 20360
rect 19706 20304 19708 20324
rect 19708 20304 19760 20324
rect 19760 20304 19762 20324
rect 19614 20168 19670 20224
rect 18878 17448 18934 17504
rect 20166 20168 20222 20224
rect 19798 18536 19854 18592
rect 19338 18028 19340 18048
rect 19340 18028 19392 18048
rect 19392 18028 19394 18048
rect 19338 17992 19394 18028
rect 19246 17584 19302 17640
rect 19154 15680 19210 15736
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 19154 15272 19210 15328
rect 19798 17992 19854 18048
rect 19706 17040 19762 17096
rect 18786 13504 18842 13560
rect 18694 12552 18750 12608
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 21086 21800 21142 21856
rect 20350 19624 20406 19680
rect 20166 17992 20222 18048
rect 20902 21392 20958 21448
rect 21086 21392 21142 21448
rect 21178 21256 21234 21312
rect 21086 20304 21142 20360
rect 20258 17604 20314 17640
rect 20258 17584 20260 17604
rect 20260 17584 20312 17604
rect 20312 17584 20314 17604
rect 19982 15136 20038 15192
rect 20074 14320 20130 14376
rect 18510 8200 18566 8256
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19890 12824 19946 12880
rect 21086 17992 21142 18048
rect 20718 16904 20774 16960
rect 20718 16496 20774 16552
rect 20350 14320 20406 14376
rect 20258 14048 20314 14104
rect 20994 17040 21050 17096
rect 20902 16496 20958 16552
rect 21454 17856 21510 17912
rect 21454 17040 21510 17096
rect 21638 20712 21694 20768
rect 21914 20052 21970 20088
rect 21914 20032 21916 20052
rect 21916 20032 21968 20052
rect 21968 20032 21970 20052
rect 21730 19080 21786 19136
rect 21638 17604 21694 17640
rect 21638 17584 21640 17604
rect 21640 17584 21692 17604
rect 21692 17584 21694 17604
rect 21822 15952 21878 16008
rect 21178 14864 21234 14920
rect 20810 11736 20866 11792
rect 21914 10512 21970 10568
rect 23110 26560 23166 26616
rect 22466 23568 22522 23624
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 23386 24384 23442 24440
rect 22466 19508 22522 19544
rect 22466 19488 22468 19508
rect 22468 19488 22520 19508
rect 22520 19488 22522 19508
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23202 21800 23258 21856
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23478 22480 23534 22536
rect 23846 23060 23848 23080
rect 23848 23060 23900 23080
rect 23900 23060 23902 23080
rect 23846 23024 23902 23060
rect 23294 20712 23350 20768
rect 23662 21120 23718 21176
rect 24030 23024 24086 23080
rect 25134 26288 25190 26344
rect 24674 22616 24730 22672
rect 23570 20596 23626 20632
rect 23570 20576 23572 20596
rect 23572 20576 23624 20596
rect 23624 20576 23626 20596
rect 23570 20304 23626 20360
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22282 13504 22338 13560
rect 22558 15000 22614 15056
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22466 11056 22522 11112
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 23662 17176 23718 17232
rect 23938 17992 23994 18048
rect 24030 17040 24086 17096
rect 23662 15272 23718 15328
rect 23386 13524 23442 13560
rect 23386 13504 23388 13524
rect 23388 13504 23440 13524
rect 23440 13504 23442 13524
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 23754 13504 23810 13560
rect 24122 14068 24178 14104
rect 24122 14048 24124 14068
rect 24124 14048 24176 14068
rect 24176 14048 24178 14068
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 24214 12688 24270 12744
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22374 7792 22430 7848
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 25134 22924 25136 22944
rect 25136 22924 25188 22944
rect 25188 22924 25190 22944
rect 25134 22888 25190 22924
rect 25410 23432 25466 23488
rect 24950 21836 24952 21856
rect 24952 21836 25004 21856
rect 25004 21836 25006 21856
rect 24950 21800 25006 21836
rect 25226 21256 25282 21312
rect 25870 24656 25926 24712
rect 24766 17876 24822 17912
rect 24766 17856 24768 17876
rect 24768 17856 24820 17876
rect 24820 17856 24822 17876
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 24950 14456 25006 14512
rect 26330 24384 26386 24440
rect 26698 24656 26754 24712
rect 26882 24384 26938 24440
rect 26882 23976 26938 24032
rect 26698 23704 26754 23760
rect 26974 23704 27030 23760
rect 26146 22344 26202 22400
rect 25962 20052 26018 20088
rect 25962 20032 25964 20052
rect 25964 20032 26016 20052
rect 26016 20032 26018 20052
rect 27066 23296 27122 23352
rect 26606 21800 26662 21856
rect 26238 19508 26294 19544
rect 26238 19488 26240 19508
rect 26240 19488 26292 19508
rect 26292 19488 26294 19508
rect 26330 19216 26386 19272
rect 25870 17040 25926 17096
rect 25594 15136 25650 15192
rect 25502 11736 25558 11792
rect 24306 9016 24362 9072
rect 24766 7928 24822 7984
rect 22742 7112 22798 7168
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 26238 15408 26294 15464
rect 25134 7248 25190 7304
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 27342 24928 27398 24984
rect 27986 25200 28042 25256
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27710 22924 27712 22944
rect 27712 22924 27764 22944
rect 27764 22924 27766 22944
rect 27710 22888 27766 22924
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 29458 24792 29514 24848
rect 28998 24248 29054 24304
rect 29182 23976 29238 24032
rect 29366 23840 29422 23896
rect 28722 23160 28778 23216
rect 28630 22888 28686 22944
rect 27434 21664 27490 21720
rect 27710 21800 27766 21856
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 28814 22616 28870 22672
rect 28538 21528 28594 21584
rect 27710 20848 27766 20904
rect 28538 21120 28594 21176
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27802 19624 27858 19680
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27618 19488 27674 19544
rect 26882 19080 26938 19136
rect 26882 18536 26938 18592
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 28814 20848 28870 20904
rect 28630 18944 28686 19000
rect 28814 19216 28870 19272
rect 28354 17720 28410 17776
rect 28538 17720 28594 17776
rect 28354 17448 28410 17504
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 28538 17040 28594 17096
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27618 15136 27674 15192
rect 28998 16632 29054 16688
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 26882 13640 26938 13696
rect 26882 13096 26938 13152
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 29458 22752 29514 22808
rect 30930 26560 30986 26616
rect 30562 22480 30618 22536
rect 30378 21936 30434 21992
rect 30378 21256 30434 21312
rect 32126 26424 32182 26480
rect 31390 23568 31446 23624
rect 31850 23976 31906 24032
rect 30838 22072 30894 22128
rect 31666 22616 31722 22672
rect 30102 17992 30158 18048
rect 30194 17856 30250 17912
rect 30194 17176 30250 17232
rect 29642 15544 29698 15600
rect 29550 12144 29606 12200
rect 31942 21956 31998 21992
rect 31942 21936 31944 21956
rect 31944 21936 31996 21956
rect 31996 21936 31998 21956
rect 32310 23024 32366 23080
rect 32310 21548 32366 21584
rect 32310 21528 32312 21548
rect 32312 21528 32364 21548
rect 32364 21528 32366 21548
rect 31666 20032 31722 20088
rect 30654 16496 30710 16552
rect 30378 16088 30434 16144
rect 30010 11600 30066 11656
rect 31574 18808 31630 18864
rect 31758 13640 31814 13696
rect 32126 19080 32182 19136
rect 32034 17584 32090 17640
rect 32586 23432 32642 23488
rect 32862 24928 32918 24984
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32862 23860 32918 23896
rect 32862 23840 32864 23860
rect 32864 23840 32916 23860
rect 32916 23840 32918 23860
rect 33046 23704 33102 23760
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32770 22344 32826 22400
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32310 20168 32366 20224
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32862 21004 32918 21040
rect 33598 26288 33654 26344
rect 33598 22752 33654 22808
rect 33414 21684 33470 21720
rect 33414 21664 33416 21684
rect 33416 21664 33468 21684
rect 33468 21664 33470 21684
rect 32862 20984 32864 21004
rect 32864 20984 32916 21004
rect 32916 20984 32918 21004
rect 32402 19896 32458 19952
rect 32770 20440 32826 20496
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 33874 21800 33930 21856
rect 34334 24656 34390 24712
rect 34794 25880 34850 25936
rect 34886 24248 34942 24304
rect 35070 23160 35126 23216
rect 35806 25200 35862 25256
rect 35990 25472 36046 25528
rect 35530 22888 35586 22944
rect 34334 21564 34336 21584
rect 34336 21564 34388 21584
rect 34388 21564 34390 21584
rect 34334 21528 34390 21564
rect 33138 19760 33194 19816
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32678 17448 32734 17504
rect 32586 15952 32642 16008
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32862 13776 32918 13832
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 34334 20304 34390 20360
rect 33782 17720 33838 17776
rect 35346 20848 35402 20904
rect 35530 20848 35586 20904
rect 34702 14320 34758 14376
rect 33690 13912 33746 13968
rect 35070 9968 35126 10024
rect 35254 18128 35310 18184
rect 35898 21392 35954 21448
rect 35162 9424 35218 9480
rect 37002 25608 37058 25664
rect 36726 24112 36782 24168
rect 37462 25336 37518 25392
rect 37278 22480 37334 22536
rect 35990 12280 36046 12336
rect 36634 19352 36690 19408
rect 36542 9560 36598 9616
rect 36450 8880 36506 8936
rect 36726 8336 36782 8392
rect 38750 26152 38806 26208
rect 38474 25744 38530 25800
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 39118 25064 39174 25120
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 38934 19216 38990 19272
rect 37830 18672 37886 18728
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37646 13368 37702 13424
rect 37094 13232 37150 13288
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 45834 24792 45890 24848
rect 45466 23024 45522 23080
rect 46202 23704 46258 23760
rect 46846 21936 46902 21992
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 41510 12824 41566 12880
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 49146 20984 49202 21040
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 37002 7384 37058 7440
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 33322 6704 33378 6760
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 23105 26618 23171 26621
rect 30925 26618 30991 26621
rect 23105 26616 30991 26618
rect 23105 26560 23110 26616
rect 23166 26560 30930 26616
rect 30986 26560 30991 26616
rect 23105 26558 30991 26560
rect 23105 26555 23171 26558
rect 30925 26555 30991 26558
rect 19241 26482 19307 26485
rect 32121 26482 32187 26485
rect 19241 26480 32187 26482
rect 19241 26424 19246 26480
rect 19302 26424 32126 26480
rect 32182 26424 32187 26480
rect 19241 26422 32187 26424
rect 19241 26419 19307 26422
rect 32121 26419 32187 26422
rect 12566 26284 12572 26348
rect 12636 26346 12642 26348
rect 17953 26346 18019 26349
rect 12636 26344 18019 26346
rect 12636 26288 17958 26344
rect 18014 26288 18019 26344
rect 12636 26286 18019 26288
rect 12636 26284 12642 26286
rect 17953 26283 18019 26286
rect 25129 26346 25195 26349
rect 33593 26346 33659 26349
rect 25129 26344 33659 26346
rect 25129 26288 25134 26344
rect 25190 26288 33598 26344
rect 33654 26288 33659 26344
rect 25129 26286 33659 26288
rect 25129 26283 25195 26286
rect 33593 26283 33659 26286
rect 15561 26210 15627 26213
rect 38745 26210 38811 26213
rect 15561 26208 38811 26210
rect 15561 26152 15566 26208
rect 15622 26152 38750 26208
rect 38806 26152 38811 26208
rect 15561 26150 38811 26152
rect 15561 26147 15627 26150
rect 38745 26147 38811 26150
rect 13629 26074 13695 26077
rect 33358 26074 33364 26076
rect 13629 26072 33364 26074
rect 13629 26016 13634 26072
rect 13690 26016 33364 26072
rect 13629 26014 33364 26016
rect 13629 26011 13695 26014
rect 33358 26012 33364 26014
rect 33428 26012 33434 26076
rect 12750 25876 12756 25940
rect 12820 25938 12826 25940
rect 16757 25938 16823 25941
rect 12820 25936 16823 25938
rect 12820 25880 16762 25936
rect 16818 25880 16823 25936
rect 12820 25878 16823 25880
rect 12820 25876 12826 25878
rect 16757 25875 16823 25878
rect 17953 25938 18019 25941
rect 34789 25938 34855 25941
rect 17953 25936 34855 25938
rect 17953 25880 17958 25936
rect 18014 25880 34794 25936
rect 34850 25880 34855 25936
rect 17953 25878 34855 25880
rect 17953 25875 18019 25878
rect 34789 25875 34855 25878
rect 11462 25740 11468 25804
rect 11532 25802 11538 25804
rect 38469 25802 38535 25805
rect 11532 25800 38535 25802
rect 11532 25744 38474 25800
rect 38530 25744 38535 25800
rect 11532 25742 38535 25744
rect 11532 25740 11538 25742
rect 38469 25739 38535 25742
rect 0 25666 800 25696
rect 3877 25666 3943 25669
rect 0 25664 3943 25666
rect 0 25608 3882 25664
rect 3938 25608 3943 25664
rect 0 25606 3943 25608
rect 0 25576 800 25606
rect 3877 25603 3943 25606
rect 16573 25666 16639 25669
rect 36997 25666 37063 25669
rect 16573 25664 37063 25666
rect 16573 25608 16578 25664
rect 16634 25608 37002 25664
rect 37058 25608 37063 25664
rect 16573 25606 37063 25608
rect 16573 25603 16639 25606
rect 36997 25603 37063 25606
rect 7373 25530 7439 25533
rect 16614 25530 16620 25532
rect 7373 25528 16620 25530
rect 7373 25472 7378 25528
rect 7434 25472 16620 25528
rect 7373 25470 16620 25472
rect 7373 25467 7439 25470
rect 16614 25468 16620 25470
rect 16684 25468 16690 25532
rect 16757 25530 16823 25533
rect 35985 25530 36051 25533
rect 16757 25528 36051 25530
rect 16757 25472 16762 25528
rect 16818 25472 35990 25528
rect 36046 25472 36051 25528
rect 16757 25470 36051 25472
rect 16757 25467 16823 25470
rect 35985 25467 36051 25470
rect 14406 25332 14412 25396
rect 14476 25394 14482 25396
rect 37457 25394 37523 25397
rect 14476 25392 37523 25394
rect 14476 25336 37462 25392
rect 37518 25336 37523 25392
rect 14476 25334 37523 25336
rect 14476 25332 14482 25334
rect 37457 25331 37523 25334
rect 0 25258 800 25288
rect 3141 25258 3207 25261
rect 0 25256 3207 25258
rect 0 25200 3146 25256
rect 3202 25200 3207 25256
rect 0 25198 3207 25200
rect 0 25168 800 25198
rect 3141 25195 3207 25198
rect 9581 25258 9647 25261
rect 24894 25258 24900 25260
rect 9581 25256 24900 25258
rect 9581 25200 9586 25256
rect 9642 25200 24900 25256
rect 9581 25198 24900 25200
rect 9581 25195 9647 25198
rect 24894 25196 24900 25198
rect 24964 25196 24970 25260
rect 27981 25258 28047 25261
rect 35801 25258 35867 25261
rect 27981 25256 35867 25258
rect 27981 25200 27986 25256
rect 28042 25200 35806 25256
rect 35862 25200 35867 25256
rect 27981 25198 35867 25200
rect 27981 25195 28047 25198
rect 35801 25195 35867 25198
rect 14222 25060 14228 25124
rect 14292 25122 14298 25124
rect 39113 25122 39179 25125
rect 14292 25120 39179 25122
rect 14292 25064 39118 25120
rect 39174 25064 39179 25120
rect 14292 25062 39179 25064
rect 14292 25060 14298 25062
rect 39113 25059 39179 25062
rect 6453 24986 6519 24989
rect 20069 24986 20135 24989
rect 6453 24984 20135 24986
rect 6453 24928 6458 24984
rect 6514 24928 20074 24984
rect 20130 24928 20135 24984
rect 6453 24926 20135 24928
rect 6453 24923 6519 24926
rect 20069 24923 20135 24926
rect 27337 24986 27403 24989
rect 32857 24986 32923 24989
rect 27337 24984 32923 24986
rect 27337 24928 27342 24984
rect 27398 24928 32862 24984
rect 32918 24928 32923 24984
rect 27337 24926 32923 24928
rect 27337 24923 27403 24926
rect 32857 24923 32923 24926
rect 0 24850 800 24880
rect 3693 24850 3759 24853
rect 0 24848 3759 24850
rect 0 24792 3698 24848
rect 3754 24792 3759 24848
rect 0 24790 3759 24792
rect 0 24760 800 24790
rect 3693 24787 3759 24790
rect 4245 24850 4311 24853
rect 14825 24850 14891 24853
rect 4245 24848 14891 24850
rect 4245 24792 4250 24848
rect 4306 24792 14830 24848
rect 14886 24792 14891 24848
rect 4245 24790 14891 24792
rect 4245 24787 4311 24790
rect 14825 24787 14891 24790
rect 17217 24850 17283 24853
rect 29453 24850 29519 24853
rect 17217 24848 29519 24850
rect 17217 24792 17222 24848
rect 17278 24792 29458 24848
rect 29514 24792 29519 24848
rect 17217 24790 29519 24792
rect 17217 24787 17283 24790
rect 29453 24787 29519 24790
rect 45829 24850 45895 24853
rect 50200 24850 51000 24880
rect 45829 24848 51000 24850
rect 45829 24792 45834 24848
rect 45890 24792 51000 24848
rect 45829 24790 51000 24792
rect 45829 24787 45895 24790
rect 50200 24760 51000 24790
rect 3969 24714 4035 24717
rect 13721 24714 13787 24717
rect 25865 24714 25931 24717
rect 3969 24712 13554 24714
rect 3969 24656 3974 24712
rect 4030 24656 13554 24712
rect 3969 24654 13554 24656
rect 3969 24651 4035 24654
rect 13494 24578 13554 24654
rect 13721 24712 25931 24714
rect 13721 24656 13726 24712
rect 13782 24656 25870 24712
rect 25926 24656 25931 24712
rect 13721 24654 25931 24656
rect 13721 24651 13787 24654
rect 25865 24651 25931 24654
rect 26693 24714 26759 24717
rect 34329 24714 34395 24717
rect 26693 24712 34395 24714
rect 26693 24656 26698 24712
rect 26754 24656 34334 24712
rect 34390 24656 34395 24712
rect 26693 24654 34395 24656
rect 26693 24651 26759 24654
rect 34329 24651 34395 24654
rect 14549 24578 14615 24581
rect 13494 24576 14615 24578
rect 13494 24520 14554 24576
rect 14610 24520 14615 24576
rect 13494 24518 14615 24520
rect 14549 24515 14615 24518
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 12065 24442 12131 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 11838 24440 12131 24442
rect 11838 24384 12070 24440
rect 12126 24384 12131 24440
rect 11838 24382 12131 24384
rect 1577 24306 1643 24309
rect 11838 24306 11898 24382
rect 12065 24379 12131 24382
rect 15694 24380 15700 24444
rect 15764 24442 15770 24444
rect 16021 24442 16087 24445
rect 18873 24442 18939 24445
rect 15764 24440 18939 24442
rect 15764 24384 16026 24440
rect 16082 24384 18878 24440
rect 18934 24384 18939 24440
rect 15764 24382 18939 24384
rect 15764 24380 15770 24382
rect 16021 24379 16087 24382
rect 18873 24379 18939 24382
rect 23381 24442 23447 24445
rect 26325 24442 26391 24445
rect 23381 24440 26391 24442
rect 23381 24384 23386 24440
rect 23442 24384 26330 24440
rect 26386 24384 26391 24440
rect 23381 24382 26391 24384
rect 23381 24379 23447 24382
rect 26325 24379 26391 24382
rect 26877 24442 26943 24445
rect 26877 24440 31770 24442
rect 26877 24384 26882 24440
rect 26938 24384 31770 24440
rect 26877 24382 31770 24384
rect 26877 24379 26943 24382
rect 1577 24304 11898 24306
rect 1577 24248 1582 24304
rect 1638 24248 11898 24304
rect 1577 24246 11898 24248
rect 11973 24306 12039 24309
rect 28993 24306 29059 24309
rect 11973 24304 29059 24306
rect 11973 24248 11978 24304
rect 12034 24248 28998 24304
rect 29054 24248 29059 24304
rect 11973 24246 29059 24248
rect 31710 24306 31770 24382
rect 34881 24306 34947 24309
rect 31710 24304 34947 24306
rect 31710 24248 34886 24304
rect 34942 24248 34947 24304
rect 31710 24246 34947 24248
rect 1577 24243 1643 24246
rect 11973 24243 12039 24246
rect 28993 24243 29059 24246
rect 34881 24243 34947 24246
rect 1761 24170 1827 24173
rect 13721 24170 13787 24173
rect 1761 24168 13787 24170
rect 1761 24112 1766 24168
rect 1822 24112 13726 24168
rect 13782 24112 13787 24168
rect 1761 24110 13787 24112
rect 1761 24107 1827 24110
rect 13721 24107 13787 24110
rect 14549 24170 14615 24173
rect 36721 24170 36787 24173
rect 14549 24168 36787 24170
rect 14549 24112 14554 24168
rect 14610 24112 36726 24168
rect 36782 24112 36787 24168
rect 14549 24110 36787 24112
rect 14549 24107 14615 24110
rect 36721 24107 36787 24110
rect 0 24034 800 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 800 23974
rect 4061 23971 4127 23974
rect 21817 24034 21883 24037
rect 26877 24034 26943 24037
rect 21817 24032 26943 24034
rect 21817 23976 21822 24032
rect 21878 23976 26882 24032
rect 26938 23976 26943 24032
rect 21817 23974 26943 23976
rect 21817 23971 21883 23974
rect 26877 23971 26943 23974
rect 29177 24034 29243 24037
rect 31845 24034 31911 24037
rect 29177 24032 31911 24034
rect 29177 23976 29182 24032
rect 29238 23976 31850 24032
rect 31906 23976 31911 24032
rect 29177 23974 31911 23976
rect 29177 23971 29243 23974
rect 31845 23971 31911 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 11145 23898 11211 23901
rect 29361 23898 29427 23901
rect 32857 23898 32923 23901
rect 50200 23898 51000 23928
rect 11145 23896 17234 23898
rect 11145 23840 11150 23896
rect 11206 23840 17234 23896
rect 11145 23838 17234 23840
rect 11145 23835 11211 23838
rect 10041 23762 10107 23765
rect 13670 23762 13676 23764
rect 10041 23760 13676 23762
rect 10041 23704 10046 23760
rect 10102 23704 13676 23760
rect 10041 23702 13676 23704
rect 10041 23699 10107 23702
rect 13670 23700 13676 23702
rect 13740 23700 13746 23764
rect 14825 23762 14891 23765
rect 17174 23762 17234 23838
rect 29361 23896 32923 23898
rect 29361 23840 29366 23896
rect 29422 23840 32862 23896
rect 32918 23840 32923 23896
rect 29361 23838 32923 23840
rect 29361 23835 29427 23838
rect 32857 23835 32923 23838
rect 48454 23838 51000 23898
rect 26693 23762 26759 23765
rect 14825 23760 15394 23762
rect 14825 23704 14830 23760
rect 14886 23704 15394 23760
rect 14825 23702 15394 23704
rect 17174 23760 26759 23762
rect 17174 23704 26698 23760
rect 26754 23704 26759 23760
rect 17174 23702 26759 23704
rect 14825 23699 14891 23702
rect 0 23626 800 23656
rect 3969 23626 4035 23629
rect 0 23624 4035 23626
rect 0 23568 3974 23624
rect 4030 23568 4035 23624
rect 0 23566 4035 23568
rect 0 23536 800 23566
rect 3969 23563 4035 23566
rect 8109 23626 8175 23629
rect 15142 23626 15148 23628
rect 8109 23624 15148 23626
rect 8109 23568 8114 23624
rect 8170 23568 15148 23624
rect 8109 23566 15148 23568
rect 8109 23563 8175 23566
rect 15142 23564 15148 23566
rect 15212 23564 15218 23628
rect 15334 23626 15394 23702
rect 26693 23699 26759 23702
rect 26969 23762 27035 23765
rect 33041 23762 33107 23765
rect 26969 23760 33107 23762
rect 26969 23704 26974 23760
rect 27030 23704 33046 23760
rect 33102 23704 33107 23760
rect 26969 23702 33107 23704
rect 26969 23699 27035 23702
rect 33041 23699 33107 23702
rect 46197 23762 46263 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46197 23760 48514 23762
rect 46197 23704 46202 23760
rect 46258 23704 48514 23760
rect 46197 23702 48514 23704
rect 46197 23699 46263 23702
rect 19926 23626 19932 23628
rect 15334 23566 19932 23626
rect 19926 23564 19932 23566
rect 19996 23564 20002 23628
rect 22461 23626 22527 23629
rect 31385 23626 31451 23629
rect 22461 23624 31451 23626
rect 22461 23568 22466 23624
rect 22522 23568 31390 23624
rect 31446 23568 31451 23624
rect 22461 23566 31451 23568
rect 22461 23563 22527 23566
rect 31385 23563 31451 23566
rect 9305 23490 9371 23493
rect 15285 23492 15351 23493
rect 9622 23490 9628 23492
rect 9305 23488 9628 23490
rect 9305 23432 9310 23488
rect 9366 23432 9628 23488
rect 9305 23430 9628 23432
rect 9305 23427 9371 23430
rect 9622 23428 9628 23430
rect 9692 23428 9698 23492
rect 15285 23488 15332 23492
rect 15396 23490 15402 23492
rect 15653 23490 15719 23493
rect 19793 23490 19859 23493
rect 15285 23432 15290 23488
rect 15285 23428 15332 23432
rect 15396 23430 15442 23490
rect 15653 23488 19859 23490
rect 15653 23432 15658 23488
rect 15714 23432 19798 23488
rect 19854 23432 19859 23488
rect 15653 23430 19859 23432
rect 15396 23428 15402 23430
rect 15285 23427 15351 23428
rect 15653 23427 15719 23430
rect 19793 23427 19859 23430
rect 25405 23490 25471 23493
rect 32581 23490 32647 23493
rect 25405 23488 32647 23490
rect 25405 23432 25410 23488
rect 25466 23432 32586 23488
rect 32642 23432 32647 23488
rect 25405 23430 32647 23432
rect 25405 23427 25471 23430
rect 32581 23427 32647 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 27061 23354 27127 23357
rect 27061 23352 31770 23354
rect 27061 23296 27066 23352
rect 27122 23296 31770 23352
rect 27061 23294 31770 23296
rect 27061 23291 27127 23294
rect 0 23218 800 23248
rect 3877 23218 3943 23221
rect 0 23216 3943 23218
rect 0 23160 3882 23216
rect 3938 23160 3943 23216
rect 0 23158 3943 23160
rect 0 23128 800 23158
rect 3877 23155 3943 23158
rect 6821 23218 6887 23221
rect 14457 23218 14523 23221
rect 17953 23218 18019 23221
rect 28717 23218 28783 23221
rect 6821 23216 16314 23218
rect 6821 23160 6826 23216
rect 6882 23160 14462 23216
rect 14518 23160 16314 23216
rect 6821 23158 16314 23160
rect 6821 23155 6887 23158
rect 14457 23155 14523 23158
rect 4061 23082 4127 23085
rect 12617 23082 12683 23085
rect 13854 23082 13860 23084
rect 4061 23080 12450 23082
rect 4061 23024 4066 23080
rect 4122 23024 12450 23080
rect 4061 23022 12450 23024
rect 4061 23019 4127 23022
rect 9765 22946 9831 22949
rect 11462 22946 11468 22948
rect 9765 22944 11468 22946
rect 9765 22888 9770 22944
rect 9826 22888 11468 22944
rect 9765 22886 11468 22888
rect 9765 22883 9831 22886
rect 11462 22884 11468 22886
rect 11532 22884 11538 22948
rect 12390 22946 12450 23022
rect 12617 23080 13860 23082
rect 12617 23024 12622 23080
rect 12678 23024 13860 23080
rect 12617 23022 13860 23024
rect 12617 23019 12683 23022
rect 13854 23020 13860 23022
rect 13924 23020 13930 23084
rect 16254 23082 16314 23158
rect 17953 23216 28783 23218
rect 17953 23160 17958 23216
rect 18014 23160 28722 23216
rect 28778 23160 28783 23216
rect 17953 23158 28783 23160
rect 31710 23218 31770 23294
rect 35065 23218 35131 23221
rect 31710 23216 35131 23218
rect 31710 23160 35070 23216
rect 35126 23160 35131 23216
rect 31710 23158 35131 23160
rect 17953 23155 18019 23158
rect 28717 23155 28783 23158
rect 35065 23155 35131 23158
rect 23841 23082 23907 23085
rect 24025 23082 24091 23085
rect 32305 23082 32371 23085
rect 16254 23080 23907 23082
rect 16254 23024 23846 23080
rect 23902 23024 23907 23080
rect 16254 23022 23907 23024
rect 23841 23019 23907 23022
rect 23982 23080 32371 23082
rect 23982 23024 24030 23080
rect 24086 23024 32310 23080
rect 32366 23024 32371 23080
rect 23982 23022 32371 23024
rect 23982 23019 24091 23022
rect 32305 23019 32371 23022
rect 45461 23082 45527 23085
rect 45461 23080 48514 23082
rect 45461 23024 45466 23080
rect 45522 23024 48514 23080
rect 45461 23022 48514 23024
rect 45461 23019 45527 23022
rect 16849 22946 16915 22949
rect 12390 22944 16915 22946
rect 12390 22888 16854 22944
rect 16910 22888 16915 22944
rect 12390 22886 16915 22888
rect 16849 22883 16915 22886
rect 19149 22946 19215 22949
rect 23982 22946 24042 23019
rect 19149 22944 24042 22946
rect 19149 22888 19154 22944
rect 19210 22888 24042 22944
rect 19149 22886 24042 22888
rect 25129 22946 25195 22949
rect 27705 22946 27771 22949
rect 25129 22944 27771 22946
rect 25129 22888 25134 22944
rect 25190 22888 27710 22944
rect 27766 22888 27771 22944
rect 25129 22886 27771 22888
rect 19149 22883 19215 22886
rect 25129 22883 25195 22886
rect 27705 22883 27771 22886
rect 28625 22946 28691 22949
rect 35525 22946 35591 22949
rect 28625 22944 35591 22946
rect 28625 22888 28630 22944
rect 28686 22888 35530 22944
rect 35586 22888 35591 22944
rect 28625 22886 35591 22888
rect 48454 22946 48514 23022
rect 50200 22946 51000 22976
rect 48454 22886 51000 22946
rect 28625 22883 28691 22886
rect 35525 22883 35591 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 50200 22856 51000 22886
rect 47946 22815 48262 22816
rect 4061 22810 4127 22813
rect 0 22808 4127 22810
rect 0 22752 4066 22808
rect 4122 22752 4127 22808
rect 0 22750 4127 22752
rect 0 22720 800 22750
rect 4061 22747 4127 22750
rect 11053 22810 11119 22813
rect 11646 22810 11652 22812
rect 11053 22808 11652 22810
rect 11053 22752 11058 22808
rect 11114 22752 11652 22808
rect 11053 22750 11652 22752
rect 11053 22747 11119 22750
rect 11646 22748 11652 22750
rect 11716 22748 11722 22812
rect 11789 22810 11855 22813
rect 12566 22810 12572 22812
rect 11789 22808 12572 22810
rect 11789 22752 11794 22808
rect 11850 22752 12572 22808
rect 11789 22750 12572 22752
rect 11789 22747 11855 22750
rect 12566 22748 12572 22750
rect 12636 22748 12642 22812
rect 13169 22810 13235 22813
rect 17401 22810 17467 22813
rect 29453 22810 29519 22813
rect 33593 22810 33659 22813
rect 13169 22808 17467 22810
rect 13169 22752 13174 22808
rect 13230 22752 17406 22808
rect 17462 22752 17467 22808
rect 13169 22750 17467 22752
rect 13169 22747 13235 22750
rect 17401 22747 17467 22750
rect 22050 22750 24962 22810
rect 3550 22612 3556 22676
rect 3620 22674 3626 22676
rect 3969 22674 4035 22677
rect 3620 22672 4035 22674
rect 3620 22616 3974 22672
rect 4030 22616 4035 22672
rect 3620 22614 4035 22616
rect 3620 22612 3626 22614
rect 3969 22611 4035 22614
rect 6913 22674 6979 22677
rect 19977 22674 20043 22677
rect 6913 22672 20043 22674
rect 6913 22616 6918 22672
rect 6974 22616 19982 22672
rect 20038 22616 20043 22672
rect 6913 22614 20043 22616
rect 6913 22611 6979 22614
rect 19977 22611 20043 22614
rect 3509 22538 3575 22541
rect 2730 22536 3575 22538
rect 2730 22480 3514 22536
rect 3570 22480 3575 22536
rect 2730 22478 3575 22480
rect 0 22402 800 22432
rect 2730 22402 2790 22478
rect 3509 22475 3575 22478
rect 6453 22538 6519 22541
rect 13169 22538 13235 22541
rect 22050 22538 22110 22750
rect 24669 22676 24735 22677
rect 24669 22672 24716 22676
rect 24780 22674 24786 22676
rect 24902 22674 24962 22750
rect 29453 22808 33659 22810
rect 29453 22752 29458 22808
rect 29514 22752 33598 22808
rect 33654 22752 33659 22808
rect 29453 22750 33659 22752
rect 29453 22747 29519 22750
rect 33593 22747 33659 22750
rect 28809 22674 28875 22677
rect 31661 22674 31727 22677
rect 24669 22616 24674 22672
rect 24669 22612 24716 22616
rect 24780 22614 24826 22674
rect 24902 22672 28875 22674
rect 24902 22616 28814 22672
rect 28870 22616 28875 22672
rect 24902 22614 28875 22616
rect 24780 22612 24786 22614
rect 24669 22611 24735 22612
rect 28809 22611 28875 22614
rect 30422 22672 31727 22674
rect 30422 22616 31666 22672
rect 31722 22616 31727 22672
rect 30422 22614 31727 22616
rect 6453 22536 13235 22538
rect 6453 22480 6458 22536
rect 6514 22480 13174 22536
rect 13230 22480 13235 22536
rect 6453 22478 13235 22480
rect 6453 22475 6519 22478
rect 13169 22475 13235 22478
rect 13356 22478 22110 22538
rect 23473 22538 23539 22541
rect 30422 22538 30482 22614
rect 31661 22611 31727 22614
rect 23473 22536 30482 22538
rect 23473 22480 23478 22536
rect 23534 22480 30482 22536
rect 23473 22478 30482 22480
rect 30557 22538 30623 22541
rect 37273 22538 37339 22541
rect 30557 22536 37339 22538
rect 30557 22480 30562 22536
rect 30618 22480 37278 22536
rect 37334 22480 37339 22536
rect 30557 22478 37339 22480
rect 0 22342 2790 22402
rect 4613 22404 4679 22405
rect 7373 22404 7439 22405
rect 4613 22400 4660 22404
rect 4724 22402 4730 22404
rect 4613 22344 4618 22400
rect 0 22312 800 22342
rect 4613 22340 4660 22344
rect 4724 22342 4770 22402
rect 7373 22400 7420 22404
rect 7484 22402 7490 22404
rect 7373 22344 7378 22400
rect 4724 22340 4730 22342
rect 7373 22340 7420 22344
rect 7484 22342 7530 22402
rect 7484 22340 7490 22342
rect 4613 22339 4679 22340
rect 7373 22339 7439 22340
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 9489 22266 9555 22269
rect 11053 22266 11119 22269
rect 9489 22264 11119 22266
rect 9489 22208 9494 22264
rect 9550 22208 11058 22264
rect 11114 22208 11119 22264
rect 9489 22206 11119 22208
rect 9489 22203 9555 22206
rect 11053 22203 11119 22206
rect 9305 22130 9371 22133
rect 13356 22130 13416 22478
rect 23473 22475 23539 22478
rect 30557 22475 30623 22478
rect 37273 22475 37339 22478
rect 26141 22402 26207 22405
rect 32765 22402 32831 22405
rect 26141 22400 32831 22402
rect 26141 22344 26146 22400
rect 26202 22344 32770 22400
rect 32826 22344 32831 22400
rect 26141 22342 32831 22344
rect 26141 22339 26207 22342
rect 32765 22339 32831 22342
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 19609 22268 19675 22269
rect 19558 22266 19564 22268
rect 19518 22206 19564 22266
rect 19628 22264 19675 22268
rect 19670 22208 19675 22264
rect 19558 22204 19564 22206
rect 19628 22204 19675 22208
rect 19609 22203 19675 22204
rect 9305 22128 13416 22130
rect 9305 22072 9310 22128
rect 9366 22072 13416 22128
rect 9305 22070 13416 22072
rect 13813 22130 13879 22133
rect 30833 22130 30899 22133
rect 13813 22128 30899 22130
rect 13813 22072 13818 22128
rect 13874 22072 30838 22128
rect 30894 22072 30899 22128
rect 13813 22070 30899 22072
rect 9305 22067 9371 22070
rect 13813 22067 13879 22070
rect 30833 22067 30899 22070
rect 0 21994 800 22024
rect 3693 21994 3759 21997
rect 0 21992 3759 21994
rect 0 21936 3698 21992
rect 3754 21936 3759 21992
rect 0 21934 3759 21936
rect 0 21904 800 21934
rect 3693 21931 3759 21934
rect 5993 21994 6059 21997
rect 10685 21994 10751 21997
rect 14222 21994 14228 21996
rect 5993 21992 10610 21994
rect 5993 21936 5998 21992
rect 6054 21936 10610 21992
rect 5993 21934 10610 21936
rect 5993 21931 6059 21934
rect 2630 21796 2636 21860
rect 2700 21858 2706 21860
rect 5625 21858 5691 21861
rect 2700 21856 5691 21858
rect 2700 21800 5630 21856
rect 5686 21800 5691 21856
rect 2700 21798 5691 21800
rect 10550 21858 10610 21934
rect 10685 21992 14228 21994
rect 10685 21936 10690 21992
rect 10746 21936 14228 21992
rect 10685 21934 14228 21936
rect 10685 21931 10751 21934
rect 14222 21932 14228 21934
rect 14292 21932 14298 21996
rect 18873 21994 18939 21997
rect 30373 21994 30439 21997
rect 31937 21994 32003 21997
rect 15702 21992 28458 21994
rect 15702 21936 18878 21992
rect 18934 21936 28458 21992
rect 15702 21934 28458 21936
rect 11697 21858 11763 21861
rect 10550 21856 11763 21858
rect 10550 21800 11702 21856
rect 11758 21800 11763 21856
rect 10550 21798 11763 21800
rect 2700 21796 2706 21798
rect 5625 21795 5691 21798
rect 11697 21795 11763 21798
rect 13353 21858 13419 21861
rect 15702 21858 15762 21934
rect 18873 21931 18939 21934
rect 13353 21856 15762 21858
rect 13353 21800 13358 21856
rect 13414 21800 15762 21856
rect 13353 21798 15762 21800
rect 18413 21858 18479 21861
rect 21081 21858 21147 21861
rect 18413 21856 21147 21858
rect 18413 21800 18418 21856
rect 18474 21800 21086 21856
rect 21142 21800 21147 21856
rect 18413 21798 21147 21800
rect 13353 21795 13419 21798
rect 18413 21795 18479 21798
rect 21081 21795 21147 21798
rect 23197 21858 23263 21861
rect 24945 21858 25011 21861
rect 26601 21858 26667 21861
rect 27705 21858 27771 21861
rect 23197 21856 27771 21858
rect 23197 21800 23202 21856
rect 23258 21800 24950 21856
rect 25006 21800 26606 21856
rect 26662 21800 27710 21856
rect 27766 21800 27771 21856
rect 23197 21798 27771 21800
rect 28398 21858 28458 21934
rect 30373 21992 32003 21994
rect 30373 21936 30378 21992
rect 30434 21936 31942 21992
rect 31998 21936 32003 21992
rect 30373 21934 32003 21936
rect 30373 21931 30439 21934
rect 31937 21931 32003 21934
rect 46841 21994 46907 21997
rect 50200 21994 51000 22024
rect 46841 21992 51000 21994
rect 46841 21936 46846 21992
rect 46902 21936 51000 21992
rect 46841 21934 51000 21936
rect 46841 21931 46907 21934
rect 50200 21904 51000 21934
rect 33869 21858 33935 21861
rect 28398 21856 33935 21858
rect 28398 21800 33874 21856
rect 33930 21800 33935 21856
rect 28398 21798 33935 21800
rect 23197 21795 23263 21798
rect 24945 21795 25011 21798
rect 26601 21795 26667 21798
rect 27705 21795 27771 21798
rect 33869 21795 33935 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 2446 21660 2452 21724
rect 2516 21722 2522 21724
rect 3785 21722 3851 21725
rect 2516 21720 3851 21722
rect 2516 21664 3790 21720
rect 3846 21664 3851 21720
rect 2516 21662 3851 21664
rect 2516 21660 2522 21662
rect 3785 21659 3851 21662
rect 10501 21722 10567 21725
rect 11053 21722 11119 21725
rect 10501 21720 11119 21722
rect 10501 21664 10506 21720
rect 10562 21664 11058 21720
rect 11114 21664 11119 21720
rect 10501 21662 11119 21664
rect 10501 21659 10567 21662
rect 11053 21659 11119 21662
rect 13077 21722 13143 21725
rect 17125 21722 17191 21725
rect 13077 21720 17191 21722
rect 13077 21664 13082 21720
rect 13138 21664 17130 21720
rect 17186 21664 17191 21720
rect 13077 21662 17191 21664
rect 13077 21659 13143 21662
rect 17125 21659 17191 21662
rect 19517 21722 19583 21725
rect 27429 21722 27495 21725
rect 33409 21724 33475 21725
rect 19517 21720 27495 21722
rect 19517 21664 19522 21720
rect 19578 21664 27434 21720
rect 27490 21664 27495 21720
rect 19517 21662 27495 21664
rect 19517 21659 19583 21662
rect 27429 21659 27495 21662
rect 28398 21662 33242 21722
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 3417 21586 3483 21589
rect 12341 21586 12407 21589
rect 3417 21584 12407 21586
rect 3417 21528 3422 21584
rect 3478 21528 12346 21584
rect 12402 21528 12407 21584
rect 3417 21526 12407 21528
rect 3417 21523 3483 21526
rect 12341 21523 12407 21526
rect 12525 21586 12591 21589
rect 28398 21586 28458 21662
rect 12525 21584 28458 21586
rect 12525 21528 12530 21584
rect 12586 21528 28458 21584
rect 12525 21526 28458 21528
rect 28533 21586 28599 21589
rect 32305 21586 32371 21589
rect 28533 21584 32371 21586
rect 28533 21528 28538 21584
rect 28594 21528 32310 21584
rect 32366 21528 32371 21584
rect 28533 21526 32371 21528
rect 33182 21586 33242 21662
rect 33358 21660 33364 21724
rect 33428 21722 33475 21724
rect 33428 21720 33520 21722
rect 33470 21664 33520 21720
rect 33428 21662 33520 21664
rect 33428 21660 33475 21662
rect 33409 21659 33475 21660
rect 34329 21586 34395 21589
rect 33182 21584 34395 21586
rect 33182 21528 34334 21584
rect 34390 21528 34395 21584
rect 33182 21526 34395 21528
rect 12525 21523 12591 21526
rect 28533 21523 28599 21526
rect 32305 21523 32371 21526
rect 34329 21523 34395 21526
rect 5165 21450 5231 21453
rect 7925 21450 7991 21453
rect 5165 21448 7991 21450
rect 5165 21392 5170 21448
rect 5226 21392 7930 21448
rect 7986 21392 7991 21448
rect 5165 21390 7991 21392
rect 5165 21387 5231 21390
rect 7925 21387 7991 21390
rect 10726 21388 10732 21452
rect 10796 21450 10802 21452
rect 10961 21450 11027 21453
rect 14181 21450 14247 21453
rect 10796 21448 12450 21450
rect 10796 21392 10966 21448
rect 11022 21392 12450 21448
rect 10796 21390 12450 21392
rect 10796 21388 10802 21390
rect 10961 21387 11027 21390
rect 5901 21314 5967 21317
rect 10501 21314 10567 21317
rect 11145 21316 11211 21317
rect 11094 21314 11100 21316
rect 5901 21312 10567 21314
rect 5901 21256 5906 21312
rect 5962 21256 10506 21312
rect 10562 21256 10567 21312
rect 5901 21254 10567 21256
rect 11054 21254 11100 21314
rect 11164 21312 11211 21316
rect 11206 21256 11211 21312
rect 5901 21251 5967 21254
rect 10501 21251 10567 21254
rect 11094 21252 11100 21254
rect 11164 21252 11211 21256
rect 12390 21314 12450 21390
rect 12804 21448 14247 21450
rect 12804 21392 14186 21448
rect 14242 21392 14247 21448
rect 12804 21390 14247 21392
rect 12804 21314 12864 21390
rect 14181 21387 14247 21390
rect 16941 21450 17007 21453
rect 20897 21450 20963 21453
rect 16941 21448 20963 21450
rect 16941 21392 16946 21448
rect 17002 21392 20902 21448
rect 20958 21392 20963 21448
rect 16941 21390 20963 21392
rect 16941 21387 17007 21390
rect 20897 21387 20963 21390
rect 21081 21450 21147 21453
rect 35893 21450 35959 21453
rect 21081 21448 35959 21450
rect 21081 21392 21086 21448
rect 21142 21392 35898 21448
rect 35954 21392 35959 21448
rect 21081 21390 35959 21392
rect 21081 21387 21147 21390
rect 35893 21387 35959 21390
rect 12390 21254 12864 21314
rect 13670 21252 13676 21316
rect 13740 21314 13746 21316
rect 17585 21314 17651 21317
rect 13740 21312 17651 21314
rect 13740 21256 17590 21312
rect 17646 21256 17651 21312
rect 13740 21254 17651 21256
rect 13740 21252 13746 21254
rect 11145 21251 11211 21252
rect 17585 21251 17651 21254
rect 17861 21314 17927 21317
rect 21173 21314 21239 21317
rect 17861 21312 21239 21314
rect 17861 21256 17866 21312
rect 17922 21256 21178 21312
rect 21234 21256 21239 21312
rect 17861 21254 21239 21256
rect 17861 21251 17927 21254
rect 21173 21251 21239 21254
rect 25221 21314 25287 21317
rect 30373 21314 30439 21317
rect 25221 21312 30439 21314
rect 25221 21256 25226 21312
rect 25282 21256 30378 21312
rect 30434 21256 30439 21312
rect 25221 21254 30439 21256
rect 25221 21251 25287 21254
rect 30373 21251 30439 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 5809 21178 5875 21181
rect 12801 21178 12867 21181
rect 5809 21176 12867 21178
rect 5809 21120 5814 21176
rect 5870 21120 12806 21176
rect 12862 21120 12867 21176
rect 5809 21118 12867 21120
rect 5809 21115 5875 21118
rect 12801 21115 12867 21118
rect 13445 21178 13511 21181
rect 19742 21178 19748 21180
rect 13445 21176 19748 21178
rect 13445 21120 13450 21176
rect 13506 21120 19748 21176
rect 13445 21118 19748 21120
rect 13445 21115 13511 21118
rect 19742 21116 19748 21118
rect 19812 21116 19818 21180
rect 23657 21178 23723 21181
rect 28533 21178 28599 21181
rect 23657 21176 28599 21178
rect 23657 21120 23662 21176
rect 23718 21120 28538 21176
rect 28594 21120 28599 21176
rect 23657 21118 28599 21120
rect 23657 21115 23723 21118
rect 28533 21115 28599 21118
rect 6678 20980 6684 21044
rect 6748 21042 6754 21044
rect 8109 21042 8175 21045
rect 6748 21040 8175 21042
rect 6748 20984 8114 21040
rect 8170 20984 8175 21040
rect 6748 20982 8175 20984
rect 6748 20980 6754 20982
rect 8109 20979 8175 20982
rect 10409 21042 10475 21045
rect 10910 21042 10916 21044
rect 10409 21040 10916 21042
rect 10409 20984 10414 21040
rect 10470 20984 10916 21040
rect 10409 20982 10916 20984
rect 10409 20979 10475 20982
rect 10910 20980 10916 20982
rect 10980 20980 10986 21044
rect 14181 21042 14247 21045
rect 32857 21042 32923 21045
rect 14181 21040 32923 21042
rect 14181 20984 14186 21040
rect 14242 20984 32862 21040
rect 32918 20984 32923 21040
rect 14181 20982 32923 20984
rect 14181 20979 14247 20982
rect 32857 20979 32923 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 3601 20906 3667 20909
rect 12341 20906 12407 20909
rect 3601 20904 12407 20906
rect 3601 20848 3606 20904
rect 3662 20848 12346 20904
rect 12402 20848 12407 20904
rect 3601 20846 12407 20848
rect 3601 20843 3667 20846
rect 12341 20843 12407 20846
rect 14733 20906 14799 20909
rect 27705 20906 27771 20909
rect 14733 20904 27771 20906
rect 14733 20848 14738 20904
rect 14794 20848 27710 20904
rect 27766 20848 27771 20904
rect 14733 20846 27771 20848
rect 14733 20843 14799 20846
rect 27705 20843 27771 20846
rect 28809 20906 28875 20909
rect 35341 20906 35407 20909
rect 35525 20906 35591 20909
rect 28809 20904 35591 20906
rect 28809 20848 28814 20904
rect 28870 20848 35346 20904
rect 35402 20848 35530 20904
rect 35586 20848 35591 20904
rect 28809 20846 35591 20848
rect 28809 20843 28875 20846
rect 35341 20843 35407 20846
rect 35525 20843 35591 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 10593 20770 10659 20773
rect 14038 20770 14044 20772
rect 10593 20768 14044 20770
rect 10593 20712 10598 20768
rect 10654 20712 14044 20768
rect 10593 20710 14044 20712
rect 10593 20707 10659 20710
rect 14038 20708 14044 20710
rect 14108 20770 14114 20772
rect 14406 20770 14412 20772
rect 14108 20710 14412 20770
rect 14108 20708 14114 20710
rect 14406 20708 14412 20710
rect 14476 20708 14482 20772
rect 19425 20770 19491 20773
rect 21633 20770 21699 20773
rect 19425 20768 21699 20770
rect 19425 20712 19430 20768
rect 19486 20712 21638 20768
rect 21694 20712 21699 20768
rect 19425 20710 21699 20712
rect 19425 20707 19491 20710
rect 21633 20707 21699 20710
rect 22686 20708 22692 20772
rect 22756 20770 22762 20772
rect 23289 20770 23355 20773
rect 22756 20768 23355 20770
rect 22756 20712 23294 20768
rect 23350 20712 23355 20768
rect 22756 20710 23355 20712
rect 22756 20708 22762 20710
rect 23289 20707 23355 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 5758 20572 5764 20636
rect 5828 20634 5834 20636
rect 5901 20634 5967 20637
rect 5828 20632 5967 20634
rect 5828 20576 5906 20632
rect 5962 20576 5967 20632
rect 5828 20574 5967 20576
rect 5828 20572 5834 20574
rect 5901 20571 5967 20574
rect 9949 20634 10015 20637
rect 10358 20634 10364 20636
rect 9949 20632 10364 20634
rect 9949 20576 9954 20632
rect 10010 20576 10364 20632
rect 9949 20574 10364 20576
rect 9949 20571 10015 20574
rect 10358 20572 10364 20574
rect 10428 20572 10434 20636
rect 10501 20634 10567 20637
rect 15101 20634 15167 20637
rect 10501 20632 15167 20634
rect 10501 20576 10506 20632
rect 10562 20576 15106 20632
rect 15162 20576 15167 20632
rect 10501 20574 15167 20576
rect 10501 20571 10567 20574
rect 15101 20571 15167 20574
rect 18638 20572 18644 20636
rect 18708 20634 18714 20636
rect 18781 20634 18847 20637
rect 23565 20634 23631 20637
rect 18708 20632 23631 20634
rect 18708 20576 18786 20632
rect 18842 20576 23570 20632
rect 23626 20576 23631 20632
rect 18708 20574 23631 20576
rect 18708 20572 18714 20574
rect 18781 20571 18847 20574
rect 23565 20571 23631 20574
rect 1853 20498 1919 20501
rect 11973 20498 12039 20501
rect 1853 20496 12039 20498
rect 1853 20440 1858 20496
rect 1914 20440 11978 20496
rect 12034 20440 12039 20496
rect 1853 20438 12039 20440
rect 1853 20435 1919 20438
rect 11973 20435 12039 20438
rect 12525 20498 12591 20501
rect 19374 20498 19380 20500
rect 12525 20496 19380 20498
rect 12525 20440 12530 20496
rect 12586 20440 19380 20496
rect 12525 20438 19380 20440
rect 12525 20435 12591 20438
rect 19374 20436 19380 20438
rect 19444 20436 19450 20500
rect 32765 20498 32831 20501
rect 19566 20496 32831 20498
rect 19566 20440 32770 20496
rect 32826 20440 32831 20496
rect 19566 20438 32831 20440
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 6913 20362 6979 20365
rect 13353 20362 13419 20365
rect 6913 20360 13419 20362
rect 6913 20304 6918 20360
rect 6974 20304 13358 20360
rect 13414 20304 13419 20360
rect 6913 20302 13419 20304
rect 6913 20299 6979 20302
rect 13353 20299 13419 20302
rect 16021 20362 16087 20365
rect 19566 20362 19626 20438
rect 32765 20435 32831 20438
rect 16021 20360 19626 20362
rect 16021 20304 16026 20360
rect 16082 20304 19626 20360
rect 16021 20302 19626 20304
rect 19701 20362 19767 20365
rect 21081 20362 21147 20365
rect 23565 20362 23631 20365
rect 34329 20362 34395 20365
rect 19701 20360 21147 20362
rect 19701 20304 19706 20360
rect 19762 20304 21086 20360
rect 21142 20304 21147 20360
rect 19701 20302 21147 20304
rect 16021 20299 16087 20302
rect 19701 20299 19767 20302
rect 21081 20299 21147 20302
rect 22050 20302 23490 20362
rect 3601 20226 3667 20229
rect 12801 20226 12867 20229
rect 3601 20224 12867 20226
rect 3601 20168 3606 20224
rect 3662 20168 12806 20224
rect 12862 20168 12867 20224
rect 3601 20166 12867 20168
rect 3601 20163 3667 20166
rect 12801 20163 12867 20166
rect 17677 20226 17743 20229
rect 18689 20226 18755 20229
rect 17677 20224 18755 20226
rect 17677 20168 17682 20224
rect 17738 20168 18694 20224
rect 18750 20168 18755 20224
rect 17677 20166 18755 20168
rect 17677 20163 17743 20166
rect 18689 20163 18755 20166
rect 19609 20226 19675 20229
rect 20161 20226 20227 20229
rect 19609 20224 20227 20226
rect 19609 20168 19614 20224
rect 19670 20168 20166 20224
rect 20222 20168 20227 20224
rect 19609 20166 20227 20168
rect 19609 20163 19675 20166
rect 20161 20163 20227 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 16481 20090 16547 20093
rect 21909 20090 21975 20093
rect 22050 20090 22110 20302
rect 23430 20226 23490 20302
rect 23565 20360 34395 20362
rect 23565 20304 23570 20360
rect 23626 20304 34334 20360
rect 34390 20304 34395 20360
rect 23565 20302 34395 20304
rect 23565 20299 23631 20302
rect 34329 20299 34395 20302
rect 32305 20226 32371 20229
rect 23430 20224 32371 20226
rect 23430 20168 32310 20224
rect 32366 20168 32371 20224
rect 23430 20166 32371 20168
rect 32305 20163 32371 20166
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 16481 20088 22110 20090
rect 16481 20032 16486 20088
rect 16542 20032 21914 20088
rect 21970 20032 22110 20088
rect 16481 20030 22110 20032
rect 25957 20090 26023 20093
rect 31661 20090 31727 20093
rect 25957 20088 31727 20090
rect 25957 20032 25962 20088
rect 26018 20032 31666 20088
rect 31722 20032 31727 20088
rect 25957 20030 31727 20032
rect 16481 20027 16547 20030
rect 21909 20027 21975 20030
rect 25957 20027 26023 20030
rect 31661 20027 31727 20030
rect 0 19954 800 19984
rect 3325 19954 3391 19957
rect 8385 19954 8451 19957
rect 0 19952 3391 19954
rect 0 19896 3330 19952
rect 3386 19896 3391 19952
rect 0 19894 3391 19896
rect 0 19864 800 19894
rect 3325 19891 3391 19894
rect 7238 19952 8451 19954
rect 7238 19896 8390 19952
rect 8446 19896 8451 19952
rect 7238 19894 8451 19896
rect 1158 19756 1164 19820
rect 1228 19818 1234 19820
rect 7238 19818 7298 19894
rect 8385 19891 8451 19894
rect 9397 19954 9463 19957
rect 11513 19954 11579 19957
rect 9397 19952 11579 19954
rect 9397 19896 9402 19952
rect 9458 19896 11518 19952
rect 11574 19896 11579 19952
rect 9397 19894 11579 19896
rect 9397 19891 9463 19894
rect 11513 19891 11579 19894
rect 11973 19954 12039 19957
rect 12525 19954 12591 19957
rect 15745 19954 15811 19957
rect 11973 19952 12591 19954
rect 11973 19896 11978 19952
rect 12034 19896 12530 19952
rect 12586 19896 12591 19952
rect 11973 19894 12591 19896
rect 11973 19891 12039 19894
rect 12525 19891 12591 19894
rect 12804 19952 15811 19954
rect 12804 19896 15750 19952
rect 15806 19896 15811 19952
rect 12804 19894 15811 19896
rect 1228 19758 7298 19818
rect 7373 19818 7439 19821
rect 12341 19818 12407 19821
rect 12804 19818 12864 19894
rect 15745 19891 15811 19894
rect 17953 19954 18019 19957
rect 32397 19954 32463 19957
rect 17953 19952 32463 19954
rect 17953 19896 17958 19952
rect 18014 19896 32402 19952
rect 32458 19896 32463 19952
rect 17953 19894 32463 19896
rect 17953 19891 18019 19894
rect 32397 19891 32463 19894
rect 7373 19816 12864 19818
rect 7373 19760 7378 19816
rect 7434 19760 12346 19816
rect 12402 19760 12864 19816
rect 7373 19758 12864 19760
rect 12985 19818 13051 19821
rect 33133 19818 33199 19821
rect 12985 19816 33199 19818
rect 12985 19760 12990 19816
rect 13046 19760 33138 19816
rect 33194 19760 33199 19816
rect 12985 19758 33199 19760
rect 1228 19756 1234 19758
rect 7373 19755 7439 19758
rect 12341 19755 12407 19758
rect 12985 19755 13051 19758
rect 33133 19755 33199 19758
rect 1669 19682 1735 19685
rect 10685 19682 10751 19685
rect 12750 19682 12756 19684
rect 1669 19680 7850 19682
rect 1669 19624 1674 19680
rect 1730 19624 7850 19680
rect 1669 19622 7850 19624
rect 1669 19619 1735 19622
rect 0 19546 800 19576
rect 2957 19546 3023 19549
rect 0 19544 3023 19546
rect 0 19488 2962 19544
rect 3018 19488 3023 19544
rect 0 19486 3023 19488
rect 0 19456 800 19486
rect 2957 19483 3023 19486
rect 5574 19484 5580 19548
rect 5644 19546 5650 19548
rect 6269 19546 6335 19549
rect 5644 19544 6335 19546
rect 5644 19488 6274 19544
rect 6330 19488 6335 19544
rect 5644 19486 6335 19488
rect 5644 19484 5650 19486
rect 6269 19483 6335 19486
rect 3601 19410 3667 19413
rect 3734 19410 3740 19412
rect 3601 19408 3740 19410
rect 3601 19352 3606 19408
rect 3662 19352 3740 19408
rect 3601 19350 3740 19352
rect 3601 19347 3667 19350
rect 3734 19348 3740 19350
rect 3804 19348 3810 19412
rect 6126 19348 6132 19412
rect 6196 19410 6202 19412
rect 6545 19410 6611 19413
rect 6196 19408 6611 19410
rect 6196 19352 6550 19408
rect 6606 19352 6611 19408
rect 6196 19350 6611 19352
rect 7790 19410 7850 19622
rect 10685 19680 12756 19682
rect 10685 19624 10690 19680
rect 10746 19624 12756 19680
rect 10685 19622 12756 19624
rect 10685 19619 10751 19622
rect 12750 19620 12756 19622
rect 12820 19620 12826 19684
rect 20345 19682 20411 19685
rect 27797 19682 27863 19685
rect 20345 19680 27863 19682
rect 20345 19624 20350 19680
rect 20406 19624 27802 19680
rect 27858 19624 27863 19680
rect 20345 19622 27863 19624
rect 20345 19619 20411 19622
rect 27797 19619 27863 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 11513 19546 11579 19549
rect 13813 19546 13879 19549
rect 11513 19544 13879 19546
rect 11513 19488 11518 19544
rect 11574 19488 13818 19544
rect 13874 19488 13879 19544
rect 11513 19486 13879 19488
rect 11513 19483 11579 19486
rect 13813 19483 13879 19486
rect 22461 19548 22527 19549
rect 22461 19544 22508 19548
rect 22572 19546 22578 19548
rect 26233 19546 26299 19549
rect 27613 19546 27679 19549
rect 22461 19488 22466 19544
rect 22461 19484 22508 19488
rect 22572 19486 22618 19546
rect 26233 19544 27679 19546
rect 26233 19488 26238 19544
rect 26294 19488 27618 19544
rect 27674 19488 27679 19544
rect 26233 19486 27679 19488
rect 22572 19484 22578 19486
rect 22461 19483 22527 19484
rect 26233 19483 26299 19486
rect 27613 19483 27679 19486
rect 8293 19410 8359 19413
rect 7790 19408 8359 19410
rect 7790 19352 8298 19408
rect 8354 19352 8359 19408
rect 7790 19350 8359 19352
rect 6196 19348 6202 19350
rect 6545 19347 6611 19350
rect 8293 19347 8359 19350
rect 8702 19348 8708 19412
rect 8772 19410 8778 19412
rect 8845 19410 8911 19413
rect 11145 19410 11211 19413
rect 11278 19410 11284 19412
rect 8772 19408 8911 19410
rect 8772 19352 8850 19408
rect 8906 19352 8911 19408
rect 8772 19350 8911 19352
rect 8772 19348 8778 19350
rect 8845 19347 8911 19350
rect 9814 19350 10426 19410
rect 3325 19274 3391 19277
rect 9814 19274 9874 19350
rect 10133 19276 10199 19277
rect 10133 19274 10180 19276
rect 3325 19272 9874 19274
rect 3325 19216 3330 19272
rect 3386 19216 9874 19272
rect 3325 19214 9874 19216
rect 10088 19272 10180 19274
rect 10088 19216 10138 19272
rect 10088 19214 10180 19216
rect 3325 19211 3391 19214
rect 10133 19212 10180 19214
rect 10244 19212 10250 19276
rect 10366 19274 10426 19350
rect 11145 19408 11284 19410
rect 11145 19352 11150 19408
rect 11206 19352 11284 19408
rect 11145 19350 11284 19352
rect 11145 19347 11211 19350
rect 11278 19348 11284 19350
rect 11348 19348 11354 19412
rect 17033 19410 17099 19413
rect 17166 19410 17172 19412
rect 17033 19408 17172 19410
rect 17033 19352 17038 19408
rect 17094 19352 17172 19408
rect 17033 19350 17172 19352
rect 17033 19347 17099 19350
rect 17166 19348 17172 19350
rect 17236 19348 17242 19412
rect 18229 19410 18295 19413
rect 36629 19410 36695 19413
rect 18229 19408 36695 19410
rect 18229 19352 18234 19408
rect 18290 19352 36634 19408
rect 36690 19352 36695 19408
rect 18229 19350 36695 19352
rect 18229 19347 18295 19350
rect 36629 19347 36695 19350
rect 12157 19274 12223 19277
rect 17401 19274 17467 19277
rect 26325 19274 26391 19277
rect 10366 19272 15946 19274
rect 10366 19216 12162 19272
rect 12218 19216 15946 19272
rect 10366 19214 15946 19216
rect 10133 19211 10199 19212
rect 12157 19211 12223 19214
rect 0 19138 800 19168
rect 2681 19138 2747 19141
rect 0 19136 2747 19138
rect 0 19080 2686 19136
rect 2742 19080 2747 19136
rect 0 19078 2747 19080
rect 0 19048 800 19078
rect 2681 19075 2747 19078
rect 3601 19138 3667 19141
rect 10685 19138 10751 19141
rect 3601 19136 10751 19138
rect 3601 19080 3606 19136
rect 3662 19080 10690 19136
rect 10746 19080 10751 19136
rect 3601 19078 10751 19080
rect 3601 19075 3667 19078
rect 10685 19075 10751 19078
rect 10869 19138 10935 19141
rect 11789 19138 11855 19141
rect 10869 19136 11855 19138
rect 10869 19080 10874 19136
rect 10930 19080 11794 19136
rect 11850 19080 11855 19136
rect 10869 19078 11855 19080
rect 10869 19075 10935 19078
rect 11789 19075 11855 19078
rect 15510 19076 15516 19140
rect 15580 19138 15586 19140
rect 15653 19138 15719 19141
rect 15580 19136 15719 19138
rect 15580 19080 15658 19136
rect 15714 19080 15719 19136
rect 15580 19078 15719 19080
rect 15886 19138 15946 19214
rect 17401 19272 26391 19274
rect 17401 19216 17406 19272
rect 17462 19216 26330 19272
rect 26386 19216 26391 19272
rect 17401 19214 26391 19216
rect 17401 19211 17467 19214
rect 26325 19211 26391 19214
rect 28809 19274 28875 19277
rect 38929 19274 38995 19277
rect 28809 19272 38995 19274
rect 28809 19216 28814 19272
rect 28870 19216 38934 19272
rect 38990 19216 38995 19272
rect 28809 19214 38995 19216
rect 28809 19211 28875 19214
rect 38929 19211 38995 19214
rect 21725 19138 21791 19141
rect 15886 19136 21791 19138
rect 15886 19080 21730 19136
rect 21786 19080 21791 19136
rect 15886 19078 21791 19080
rect 15580 19076 15586 19078
rect 15653 19075 15719 19078
rect 21725 19075 21791 19078
rect 26877 19138 26943 19141
rect 32121 19138 32187 19141
rect 26877 19136 32187 19138
rect 26877 19080 26882 19136
rect 26938 19080 32126 19136
rect 32182 19080 32187 19136
rect 26877 19078 32187 19080
rect 26877 19075 26943 19078
rect 32121 19075 32187 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 4153 19002 4219 19005
rect 12341 19002 12407 19005
rect 4153 19000 12407 19002
rect 4153 18944 4158 19000
rect 4214 18944 12346 19000
rect 12402 18944 12407 19000
rect 4153 18942 12407 18944
rect 4153 18939 4219 18942
rect 12341 18939 12407 18942
rect 13905 19002 13971 19005
rect 17309 19002 17375 19005
rect 13905 19000 17375 19002
rect 13905 18944 13910 19000
rect 13966 18944 17314 19000
rect 17370 18944 17375 19000
rect 13905 18942 17375 18944
rect 13905 18939 13971 18942
rect 17309 18939 17375 18942
rect 24894 18940 24900 19004
rect 24964 19002 24970 19004
rect 28625 19002 28691 19005
rect 24964 19000 28691 19002
rect 24964 18944 28630 19000
rect 28686 18944 28691 19000
rect 24964 18942 28691 18944
rect 24964 18940 24970 18942
rect 28625 18939 28691 18942
rect 2589 18866 2655 18869
rect 5901 18866 5967 18869
rect 2589 18864 5967 18866
rect 2589 18808 2594 18864
rect 2650 18808 5906 18864
rect 5962 18808 5967 18864
rect 2589 18806 5967 18808
rect 2589 18803 2655 18806
rect 5901 18803 5967 18806
rect 9581 18866 9647 18869
rect 11605 18866 11671 18869
rect 9581 18864 11671 18866
rect 9581 18808 9586 18864
rect 9642 18808 11610 18864
rect 11666 18808 11671 18864
rect 9581 18806 11671 18808
rect 12344 18866 12404 18939
rect 14825 18866 14891 18869
rect 12344 18864 14891 18866
rect 12344 18808 14830 18864
rect 14886 18808 14891 18864
rect 12344 18806 14891 18808
rect 9581 18803 9647 18806
rect 11605 18803 11671 18806
rect 14825 18803 14891 18806
rect 15469 18866 15535 18869
rect 31569 18866 31635 18869
rect 15469 18864 31635 18866
rect 15469 18808 15474 18864
rect 15530 18808 31574 18864
rect 31630 18808 31635 18864
rect 15469 18806 31635 18808
rect 15469 18803 15535 18806
rect 31569 18803 31635 18806
rect 0 18730 800 18760
rect 2865 18730 2931 18733
rect 8293 18732 8359 18733
rect 8293 18730 8340 18732
rect 0 18728 2931 18730
rect 0 18672 2870 18728
rect 2926 18672 2931 18728
rect 0 18670 2931 18672
rect 8248 18728 8340 18730
rect 8248 18672 8298 18728
rect 8248 18670 8340 18672
rect 0 18640 800 18670
rect 2865 18667 2931 18670
rect 8293 18668 8340 18670
rect 8404 18668 8410 18732
rect 9673 18730 9739 18733
rect 10593 18730 10659 18733
rect 37825 18730 37891 18733
rect 9673 18728 10058 18730
rect 9673 18672 9678 18728
rect 9734 18672 10058 18728
rect 9673 18670 10058 18672
rect 8293 18667 8359 18668
rect 9673 18667 9739 18670
rect 1342 18532 1348 18596
rect 1412 18594 1418 18596
rect 5441 18594 5507 18597
rect 7281 18596 7347 18597
rect 1412 18592 5507 18594
rect 1412 18536 5446 18592
rect 5502 18536 5507 18592
rect 1412 18534 5507 18536
rect 1412 18532 1418 18534
rect 5441 18531 5507 18534
rect 7230 18532 7236 18596
rect 7300 18594 7347 18596
rect 9765 18596 9831 18597
rect 9765 18594 9812 18596
rect 7300 18592 7392 18594
rect 7342 18536 7392 18592
rect 7300 18534 7392 18536
rect 9720 18592 9812 18594
rect 9720 18536 9770 18592
rect 9720 18534 9812 18536
rect 7300 18532 7347 18534
rect 7281 18531 7347 18532
rect 9765 18532 9812 18534
rect 9876 18532 9882 18596
rect 9998 18594 10058 18670
rect 10593 18728 37891 18730
rect 10593 18672 10598 18728
rect 10654 18672 37830 18728
rect 37886 18672 37891 18728
rect 10593 18670 37891 18672
rect 10593 18667 10659 18670
rect 37825 18667 37891 18670
rect 9998 18534 11116 18594
rect 9765 18531 9831 18532
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 974 18396 980 18460
rect 1044 18458 1050 18460
rect 7005 18458 7071 18461
rect 1044 18456 7071 18458
rect 1044 18400 7010 18456
rect 7066 18400 7071 18456
rect 1044 18398 7071 18400
rect 11056 18458 11116 18534
rect 12014 18532 12020 18596
rect 12084 18594 12090 18596
rect 14089 18594 14155 18597
rect 12084 18592 14155 18594
rect 12084 18536 14094 18592
rect 14150 18536 14155 18592
rect 12084 18534 14155 18536
rect 12084 18532 12090 18534
rect 14089 18531 14155 18534
rect 15929 18594 15995 18597
rect 16941 18594 17007 18597
rect 15929 18592 17007 18594
rect 15929 18536 15934 18592
rect 15990 18536 16946 18592
rect 17002 18536 17007 18592
rect 15929 18534 17007 18536
rect 15929 18531 15995 18534
rect 16941 18531 17007 18534
rect 19793 18594 19859 18597
rect 26877 18594 26943 18597
rect 19793 18592 26943 18594
rect 19793 18536 19798 18592
rect 19854 18536 26882 18592
rect 26938 18536 26943 18592
rect 19793 18534 26943 18536
rect 19793 18531 19859 18534
rect 26877 18531 26943 18534
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 11605 18458 11671 18461
rect 11056 18456 11671 18458
rect 11056 18400 11610 18456
rect 11666 18400 11671 18456
rect 11056 18398 11671 18400
rect 1044 18396 1050 18398
rect 7005 18395 7071 18398
rect 11605 18395 11671 18398
rect 11789 18460 11855 18461
rect 11789 18456 11836 18460
rect 11900 18458 11906 18460
rect 12065 18458 12131 18461
rect 11900 18456 12131 18458
rect 11789 18400 11794 18456
rect 11900 18400 12070 18456
rect 12126 18400 12131 18456
rect 11789 18396 11836 18400
rect 11900 18398 12131 18400
rect 11900 18396 11906 18398
rect 11789 18395 11855 18396
rect 12065 18395 12131 18398
rect 12198 18396 12204 18460
rect 12268 18458 12274 18460
rect 13353 18458 13419 18461
rect 12268 18456 13419 18458
rect 12268 18400 13358 18456
rect 13414 18400 13419 18456
rect 12268 18398 13419 18400
rect 12268 18396 12274 18398
rect 13353 18395 13419 18398
rect 13813 18458 13879 18461
rect 17401 18458 17467 18461
rect 13813 18456 17467 18458
rect 13813 18400 13818 18456
rect 13874 18400 17406 18456
rect 17462 18400 17467 18456
rect 13813 18398 17467 18400
rect 13813 18395 13879 18398
rect 17401 18395 17467 18398
rect 0 18322 800 18352
rect 2773 18322 2839 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 0 18232 800 18262
rect 2773 18259 2839 18262
rect 8201 18322 8267 18325
rect 9990 18322 9996 18324
rect 8201 18320 9996 18322
rect 8201 18264 8206 18320
rect 8262 18264 9996 18320
rect 8201 18262 9996 18264
rect 8201 18259 8267 18262
rect 9990 18260 9996 18262
rect 10060 18322 10066 18324
rect 10685 18322 10751 18325
rect 10060 18320 10751 18322
rect 10060 18264 10690 18320
rect 10746 18264 10751 18320
rect 10060 18262 10751 18264
rect 10060 18260 10066 18262
rect 10685 18259 10751 18262
rect 11145 18322 11211 18325
rect 11513 18322 11579 18325
rect 11145 18320 11579 18322
rect 11145 18264 11150 18320
rect 11206 18264 11518 18320
rect 11574 18264 11579 18320
rect 11145 18262 11579 18264
rect 11145 18259 11211 18262
rect 11513 18259 11579 18262
rect 11789 18322 11855 18325
rect 15510 18322 15516 18324
rect 11789 18320 15516 18322
rect 11789 18264 11794 18320
rect 11850 18264 15516 18320
rect 11789 18262 15516 18264
rect 11789 18259 11855 18262
rect 15510 18260 15516 18262
rect 15580 18260 15586 18324
rect 5349 18186 5415 18189
rect 8109 18186 8175 18189
rect 8569 18188 8635 18189
rect 8518 18186 8524 18188
rect 5349 18184 8524 18186
rect 8588 18184 8635 18188
rect 5349 18128 5354 18184
rect 5410 18128 8114 18184
rect 8170 18128 8524 18184
rect 8630 18128 8635 18184
rect 5349 18126 8524 18128
rect 5349 18123 5415 18126
rect 8109 18123 8175 18126
rect 8518 18124 8524 18126
rect 8588 18124 8635 18128
rect 8569 18123 8635 18124
rect 10317 18186 10383 18189
rect 12985 18186 13051 18189
rect 16849 18186 16915 18189
rect 35249 18186 35315 18189
rect 10317 18184 16682 18186
rect 10317 18128 10322 18184
rect 10378 18128 12990 18184
rect 13046 18128 16682 18184
rect 10317 18126 16682 18128
rect 10317 18123 10383 18126
rect 12985 18123 13051 18126
rect 4102 17988 4108 18052
rect 4172 18050 4178 18052
rect 7833 18050 7899 18053
rect 4172 18048 7899 18050
rect 4172 17992 7838 18048
rect 7894 17992 7899 18048
rect 4172 17990 7899 17992
rect 4172 17988 4178 17990
rect 7833 17987 7899 17990
rect 9581 18050 9647 18053
rect 10593 18050 10659 18053
rect 9581 18048 10659 18050
rect 9581 17992 9586 18048
rect 9642 17992 10598 18048
rect 10654 17992 10659 18048
rect 9581 17990 10659 17992
rect 9581 17987 9647 17990
rect 10593 17987 10659 17990
rect 11145 18050 11211 18053
rect 12341 18050 12407 18053
rect 12801 18050 12867 18053
rect 16297 18052 16363 18053
rect 11145 18048 12867 18050
rect 11145 17992 11150 18048
rect 11206 17992 12346 18048
rect 12402 17992 12806 18048
rect 12862 17992 12867 18048
rect 11145 17990 12867 17992
rect 11145 17987 11211 17990
rect 12341 17987 12407 17990
rect 12801 17987 12867 17990
rect 16246 17988 16252 18052
rect 16316 18050 16363 18052
rect 16316 18048 16408 18050
rect 16358 17992 16408 18048
rect 16316 17990 16408 17992
rect 16316 17988 16363 17990
rect 16297 17987 16363 17988
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 4470 17852 4476 17916
rect 4540 17914 4546 17916
rect 5165 17914 5231 17917
rect 4540 17912 5231 17914
rect 4540 17856 5170 17912
rect 5226 17856 5231 17912
rect 4540 17854 5231 17856
rect 4540 17852 4546 17854
rect 5165 17851 5231 17854
rect 5993 17914 6059 17917
rect 7925 17914 7991 17917
rect 5993 17912 7991 17914
rect 5993 17856 5998 17912
rect 6054 17856 7930 17912
rect 7986 17856 7991 17912
rect 5993 17854 7991 17856
rect 5993 17851 6059 17854
rect 7925 17851 7991 17854
rect 9673 17914 9739 17917
rect 10869 17914 10935 17917
rect 9673 17912 10935 17914
rect 9673 17856 9678 17912
rect 9734 17856 10874 17912
rect 10930 17856 10935 17912
rect 9673 17854 10935 17856
rect 16622 17914 16682 18126
rect 16849 18184 35315 18186
rect 16849 18128 16854 18184
rect 16910 18128 35254 18184
rect 35310 18128 35315 18184
rect 16849 18126 35315 18128
rect 16849 18123 16915 18126
rect 35249 18123 35315 18126
rect 18413 18052 18479 18053
rect 18413 18048 18460 18052
rect 18524 18050 18530 18052
rect 19333 18050 19399 18053
rect 19793 18050 19859 18053
rect 18413 17992 18418 18048
rect 18413 17988 18460 17992
rect 18524 17990 18570 18050
rect 19333 18048 19859 18050
rect 19333 17992 19338 18048
rect 19394 17992 19798 18048
rect 19854 17992 19859 18048
rect 19333 17990 19859 17992
rect 18524 17988 18530 17990
rect 18413 17987 18479 17988
rect 19333 17987 19399 17990
rect 19793 17987 19859 17990
rect 20161 18050 20227 18053
rect 21081 18050 21147 18053
rect 20161 18048 21147 18050
rect 20161 17992 20166 18048
rect 20222 17992 21086 18048
rect 21142 17992 21147 18048
rect 20161 17990 21147 17992
rect 20161 17987 20227 17990
rect 21081 17987 21147 17990
rect 23933 18050 23999 18053
rect 30097 18050 30163 18053
rect 23933 18048 30163 18050
rect 23933 17992 23938 18048
rect 23994 17992 30102 18048
rect 30158 17992 30163 18048
rect 23933 17990 30163 17992
rect 23933 17987 23999 17990
rect 30097 17987 30163 17990
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 21449 17914 21515 17917
rect 16622 17912 21515 17914
rect 16622 17856 21454 17912
rect 21510 17856 21515 17912
rect 16622 17854 21515 17856
rect 9673 17851 9739 17854
rect 10869 17851 10935 17854
rect 21449 17851 21515 17854
rect 24761 17914 24827 17917
rect 30189 17914 30255 17917
rect 24761 17912 30255 17914
rect 24761 17856 24766 17912
rect 24822 17856 30194 17912
rect 30250 17856 30255 17912
rect 24761 17854 30255 17856
rect 24761 17851 24827 17854
rect 30189 17851 30255 17854
rect 3325 17778 3391 17781
rect 14457 17778 14523 17781
rect 3325 17776 14523 17778
rect 3325 17720 3330 17776
rect 3386 17720 14462 17776
rect 14518 17720 14523 17776
rect 3325 17718 14523 17720
rect 3325 17715 3391 17718
rect 14457 17715 14523 17718
rect 16389 17778 16455 17781
rect 28349 17778 28415 17781
rect 16389 17776 28415 17778
rect 16389 17720 16394 17776
rect 16450 17720 28354 17776
rect 28410 17720 28415 17776
rect 16389 17718 28415 17720
rect 16389 17715 16455 17718
rect 28349 17715 28415 17718
rect 28533 17778 28599 17781
rect 33777 17778 33843 17781
rect 28533 17776 33843 17778
rect 28533 17720 28538 17776
rect 28594 17720 33782 17776
rect 33838 17720 33843 17776
rect 28533 17718 33843 17720
rect 28533 17715 28599 17718
rect 33777 17715 33843 17718
rect 3918 17580 3924 17644
rect 3988 17642 3994 17644
rect 4061 17642 4127 17645
rect 3988 17640 4127 17642
rect 3988 17584 4066 17640
rect 4122 17584 4127 17640
rect 3988 17582 4127 17584
rect 3988 17580 3994 17582
rect 4061 17579 4127 17582
rect 7005 17642 7071 17645
rect 14641 17642 14707 17645
rect 7005 17640 14707 17642
rect 7005 17584 7010 17640
rect 7066 17584 14646 17640
rect 14702 17584 14707 17640
rect 7005 17582 14707 17584
rect 7005 17579 7071 17582
rect 14641 17579 14707 17582
rect 16246 17580 16252 17644
rect 16316 17642 16322 17644
rect 18229 17642 18295 17645
rect 19241 17642 19307 17645
rect 16316 17640 19307 17642
rect 16316 17584 18234 17640
rect 18290 17584 19246 17640
rect 19302 17584 19307 17640
rect 16316 17582 19307 17584
rect 16316 17580 16322 17582
rect 18229 17579 18295 17582
rect 19241 17579 19307 17582
rect 20253 17642 20319 17645
rect 21633 17642 21699 17645
rect 32029 17642 32095 17645
rect 20253 17640 21699 17642
rect 20253 17584 20258 17640
rect 20314 17584 21638 17640
rect 21694 17584 21699 17640
rect 20253 17582 21699 17584
rect 20253 17579 20319 17582
rect 21633 17579 21699 17582
rect 22050 17640 32095 17642
rect 22050 17584 32034 17640
rect 32090 17584 32095 17640
rect 22050 17582 32095 17584
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 11053 17506 11119 17509
rect 12433 17506 12499 17509
rect 11053 17504 12499 17506
rect 11053 17448 11058 17504
rect 11114 17448 12438 17504
rect 12494 17448 12499 17504
rect 11053 17446 12499 17448
rect 11053 17443 11119 17446
rect 12433 17443 12499 17446
rect 18873 17506 18939 17509
rect 22050 17506 22110 17582
rect 32029 17579 32095 17582
rect 18873 17504 22110 17506
rect 18873 17448 18878 17504
rect 18934 17448 22110 17504
rect 18873 17446 22110 17448
rect 28349 17506 28415 17509
rect 32673 17506 32739 17509
rect 28349 17504 32739 17506
rect 28349 17448 28354 17504
rect 28410 17448 32678 17504
rect 32734 17448 32739 17504
rect 28349 17446 32739 17448
rect 18873 17443 18939 17446
rect 28349 17443 28415 17446
rect 32673 17443 32739 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 9438 17308 9444 17372
rect 9508 17370 9514 17372
rect 9806 17370 9812 17372
rect 9508 17310 9812 17370
rect 9508 17308 9514 17310
rect 9806 17308 9812 17310
rect 9876 17308 9882 17372
rect 10225 17370 10291 17373
rect 15745 17370 15811 17373
rect 10225 17368 15811 17370
rect 10225 17312 10230 17368
rect 10286 17312 15750 17368
rect 15806 17312 15811 17368
rect 10225 17310 15811 17312
rect 10225 17307 10291 17310
rect 15745 17307 15811 17310
rect 1526 17172 1532 17236
rect 1596 17234 1602 17236
rect 3550 17234 3556 17236
rect 1596 17174 3556 17234
rect 1596 17172 1602 17174
rect 3550 17172 3556 17174
rect 3620 17234 3626 17236
rect 13721 17234 13787 17237
rect 3620 17232 13787 17234
rect 3620 17176 13726 17232
rect 13782 17176 13787 17232
rect 3620 17174 13787 17176
rect 3620 17172 3626 17174
rect 13721 17171 13787 17174
rect 23657 17234 23723 17237
rect 30189 17234 30255 17237
rect 23657 17232 30255 17234
rect 23657 17176 23662 17232
rect 23718 17176 30194 17232
rect 30250 17176 30255 17232
rect 23657 17174 30255 17176
rect 23657 17171 23723 17174
rect 30189 17171 30255 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 5022 17036 5028 17100
rect 5092 17098 5098 17100
rect 5625 17098 5691 17101
rect 5092 17096 13554 17098
rect 5092 17040 5630 17096
rect 5686 17040 13554 17096
rect 5092 17038 13554 17040
rect 5092 17036 5098 17038
rect 5625 17035 5691 17038
rect 7925 16962 7991 16965
rect 11789 16962 11855 16965
rect 7925 16960 11855 16962
rect 7925 16904 7930 16960
rect 7986 16904 11794 16960
rect 11850 16904 11855 16960
rect 7925 16902 11855 16904
rect 13494 16962 13554 17038
rect 14774 17036 14780 17100
rect 14844 17098 14850 17100
rect 19701 17098 19767 17101
rect 14844 17096 19767 17098
rect 14844 17040 19706 17096
rect 19762 17040 19767 17096
rect 14844 17038 19767 17040
rect 14844 17036 14850 17038
rect 19701 17035 19767 17038
rect 20989 17098 21055 17101
rect 21449 17098 21515 17101
rect 24025 17098 24091 17101
rect 20989 17096 24091 17098
rect 20989 17040 20994 17096
rect 21050 17040 21454 17096
rect 21510 17040 24030 17096
rect 24086 17040 24091 17096
rect 20989 17038 24091 17040
rect 20989 17035 21055 17038
rect 21449 17035 21515 17038
rect 24025 17035 24091 17038
rect 25865 17098 25931 17101
rect 28533 17098 28599 17101
rect 25865 17096 28599 17098
rect 25865 17040 25870 17096
rect 25926 17040 28538 17096
rect 28594 17040 28599 17096
rect 25865 17038 28599 17040
rect 25865 17035 25931 17038
rect 28533 17035 28599 17038
rect 16021 16962 16087 16965
rect 13494 16960 16087 16962
rect 13494 16904 16026 16960
rect 16082 16904 16087 16960
rect 13494 16902 16087 16904
rect 7925 16899 7991 16902
rect 11789 16899 11855 16902
rect 16021 16899 16087 16902
rect 16757 16962 16823 16965
rect 20713 16962 20779 16965
rect 16757 16960 20779 16962
rect 16757 16904 16762 16960
rect 16818 16904 20718 16960
rect 20774 16904 20779 16960
rect 16757 16902 20779 16904
rect 16757 16899 16823 16902
rect 20713 16899 20779 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 6361 16826 6427 16829
rect 8845 16826 8911 16829
rect 6361 16824 8911 16826
rect 6361 16768 6366 16824
rect 6422 16768 8850 16824
rect 8906 16768 8911 16824
rect 6361 16766 8911 16768
rect 6361 16763 6427 16766
rect 8845 16763 8911 16766
rect 9254 16764 9260 16828
rect 9324 16826 9330 16828
rect 9397 16826 9463 16829
rect 9324 16824 9463 16826
rect 9324 16768 9402 16824
rect 9458 16768 9463 16824
rect 9324 16766 9463 16768
rect 9324 16764 9330 16766
rect 9397 16763 9463 16766
rect 10593 16826 10659 16829
rect 12198 16826 12204 16828
rect 10593 16824 12204 16826
rect 10593 16768 10598 16824
rect 10654 16768 12204 16824
rect 10593 16766 12204 16768
rect 10593 16763 10659 16766
rect 12198 16764 12204 16766
rect 12268 16764 12274 16828
rect 18689 16826 18755 16829
rect 13862 16824 18755 16826
rect 13862 16768 18694 16824
rect 18750 16768 18755 16824
rect 13862 16766 18755 16768
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 3417 16690 3483 16693
rect 8109 16690 8175 16693
rect 13862 16690 13922 16766
rect 18689 16763 18755 16766
rect 3417 16688 13922 16690
rect 3417 16632 3422 16688
rect 3478 16632 8114 16688
rect 8170 16632 13922 16688
rect 3417 16630 13922 16632
rect 14089 16690 14155 16693
rect 28993 16690 29059 16693
rect 14089 16688 29059 16690
rect 14089 16632 14094 16688
rect 14150 16632 28998 16688
rect 29054 16632 29059 16688
rect 14089 16630 29059 16632
rect 3417 16627 3483 16630
rect 8109 16627 8175 16630
rect 14089 16627 14155 16630
rect 28993 16627 29059 16630
rect 5441 16554 5507 16557
rect 13813 16554 13879 16557
rect 5441 16552 13879 16554
rect 5441 16496 5446 16552
rect 5502 16496 13818 16552
rect 13874 16496 13879 16552
rect 5441 16494 13879 16496
rect 5441 16491 5507 16494
rect 13813 16491 13879 16494
rect 17309 16554 17375 16557
rect 20713 16554 20779 16557
rect 17309 16552 20779 16554
rect 17309 16496 17314 16552
rect 17370 16496 20718 16552
rect 20774 16496 20779 16552
rect 17309 16494 20779 16496
rect 17309 16491 17375 16494
rect 20713 16491 20779 16494
rect 20897 16554 20963 16557
rect 30649 16554 30715 16557
rect 20897 16552 30715 16554
rect 20897 16496 20902 16552
rect 20958 16496 30654 16552
rect 30710 16496 30715 16552
rect 20897 16494 30715 16496
rect 20897 16491 20963 16494
rect 30649 16491 30715 16494
rect 1117 16418 1183 16421
rect 7741 16418 7807 16421
rect 1117 16416 7807 16418
rect 1117 16360 1122 16416
rect 1178 16360 7746 16416
rect 7802 16360 7807 16416
rect 1117 16358 7807 16360
rect 1117 16355 1183 16358
rect 7741 16355 7807 16358
rect 9949 16418 10015 16421
rect 11789 16418 11855 16421
rect 13629 16418 13695 16421
rect 9949 16416 11668 16418
rect 9949 16360 9954 16416
rect 10010 16360 11668 16416
rect 9949 16358 11668 16360
rect 9949 16355 10015 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 5625 16282 5691 16285
rect 6085 16282 6151 16285
rect 11053 16282 11119 16285
rect 11421 16282 11487 16285
rect 5625 16280 7298 16282
rect 5625 16224 5630 16280
rect 5686 16224 6090 16280
rect 6146 16224 7298 16280
rect 5625 16222 7298 16224
rect 5625 16219 5691 16222
rect 6085 16219 6151 16222
rect 1117 16146 1183 16149
rect 7097 16146 7163 16149
rect 1117 16144 7163 16146
rect 1117 16088 1122 16144
rect 1178 16088 7102 16144
rect 7158 16088 7163 16144
rect 1117 16086 7163 16088
rect 7238 16146 7298 16222
rect 11053 16280 11487 16282
rect 11053 16224 11058 16280
rect 11114 16224 11426 16280
rect 11482 16224 11487 16280
rect 11053 16222 11487 16224
rect 11608 16282 11668 16358
rect 11789 16416 13695 16418
rect 11789 16360 11794 16416
rect 11850 16360 13634 16416
rect 13690 16360 13695 16416
rect 11789 16358 13695 16360
rect 11789 16355 11855 16358
rect 13629 16355 13695 16358
rect 13854 16356 13860 16420
rect 13924 16418 13930 16420
rect 14457 16418 14523 16421
rect 13924 16416 14523 16418
rect 13924 16360 14462 16416
rect 14518 16360 14523 16416
rect 13924 16358 14523 16360
rect 13924 16356 13930 16358
rect 14457 16355 14523 16358
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 12014 16282 12020 16284
rect 11608 16222 12020 16282
rect 11053 16219 11119 16222
rect 11421 16219 11487 16222
rect 12014 16220 12020 16222
rect 12084 16220 12090 16284
rect 12341 16282 12407 16285
rect 13813 16282 13879 16285
rect 12341 16280 13879 16282
rect 12341 16224 12346 16280
rect 12402 16224 13818 16280
rect 13874 16224 13879 16280
rect 12341 16222 13879 16224
rect 12341 16219 12407 16222
rect 13813 16219 13879 16222
rect 30373 16146 30439 16149
rect 7238 16144 30439 16146
rect 7238 16088 30378 16144
rect 30434 16088 30439 16144
rect 7238 16086 30439 16088
rect 1117 16083 1183 16086
rect 7097 16083 7163 16086
rect 30373 16083 30439 16086
rect 4153 16010 4219 16013
rect 9397 16010 9463 16013
rect 4153 16008 9463 16010
rect 4153 15952 4158 16008
rect 4214 15952 9402 16008
rect 9458 15952 9463 16008
rect 4153 15950 9463 15952
rect 4153 15947 4219 15950
rect 9397 15947 9463 15950
rect 10501 16010 10567 16013
rect 14089 16010 14155 16013
rect 21817 16010 21883 16013
rect 32581 16010 32647 16013
rect 10501 16008 13968 16010
rect 10501 15952 10506 16008
rect 10562 15952 13968 16008
rect 10501 15950 13968 15952
rect 10501 15947 10567 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 4705 15874 4771 15877
rect 5809 15874 5875 15877
rect 8477 15876 8543 15877
rect 8477 15874 8524 15876
rect 4705 15872 5875 15874
rect 4705 15816 4710 15872
rect 4766 15816 5814 15872
rect 5870 15816 5875 15872
rect 4705 15814 5875 15816
rect 8432 15872 8524 15874
rect 8432 15816 8482 15872
rect 8432 15814 8524 15816
rect 4705 15811 4771 15814
rect 5809 15811 5875 15814
rect 8477 15812 8524 15814
rect 8588 15812 8594 15876
rect 8886 15812 8892 15876
rect 8956 15874 8962 15876
rect 9581 15874 9647 15877
rect 8956 15872 9647 15874
rect 8956 15816 9586 15872
rect 9642 15816 9647 15872
rect 8956 15814 9647 15816
rect 8956 15812 8962 15814
rect 8477 15811 8543 15812
rect 9581 15811 9647 15814
rect 10961 15874 11027 15877
rect 13908 15874 13968 15950
rect 14089 16008 21883 16010
rect 14089 15952 14094 16008
rect 14150 15952 21822 16008
rect 21878 15952 21883 16008
rect 14089 15950 21883 15952
rect 14089 15947 14155 15950
rect 21817 15947 21883 15950
rect 22050 16008 32647 16010
rect 22050 15952 32586 16008
rect 32642 15952 32647 16008
rect 22050 15950 32647 15952
rect 17217 15874 17283 15877
rect 10961 15872 12864 15874
rect 10961 15816 10966 15872
rect 11022 15816 12864 15872
rect 10961 15814 12864 15816
rect 13908 15872 17283 15874
rect 13908 15816 17222 15872
rect 17278 15816 17283 15872
rect 13908 15814 17283 15816
rect 10961 15811 11027 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 5165 15738 5231 15741
rect 12433 15738 12499 15741
rect 5165 15736 12499 15738
rect 5165 15680 5170 15736
rect 5226 15680 12438 15736
rect 12494 15680 12499 15736
rect 5165 15678 12499 15680
rect 5165 15675 5231 15678
rect 12433 15675 12499 15678
rect 4429 15602 4495 15605
rect 5993 15602 6059 15605
rect 4429 15600 6059 15602
rect 4429 15544 4434 15600
rect 4490 15544 5998 15600
rect 6054 15544 6059 15600
rect 4429 15542 6059 15544
rect 4429 15539 4495 15542
rect 5993 15539 6059 15542
rect 6361 15602 6427 15605
rect 7557 15602 7623 15605
rect 12525 15602 12591 15605
rect 6361 15600 12591 15602
rect 6361 15544 6366 15600
rect 6422 15544 7562 15600
rect 7618 15544 12530 15600
rect 12586 15544 12591 15600
rect 6361 15542 12591 15544
rect 12804 15602 12864 15814
rect 17217 15811 17283 15814
rect 19374 15812 19380 15876
rect 19444 15874 19450 15876
rect 22050 15874 22110 15950
rect 32581 15947 32647 15950
rect 19444 15814 22110 15874
rect 19444 15812 19450 15814
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 14825 15738 14891 15741
rect 19149 15738 19215 15741
rect 14825 15736 19215 15738
rect 14825 15680 14830 15736
rect 14886 15680 19154 15736
rect 19210 15680 19215 15736
rect 14825 15678 19215 15680
rect 14825 15675 14891 15678
rect 19149 15675 19215 15678
rect 29637 15602 29703 15605
rect 12804 15600 29703 15602
rect 12804 15544 29642 15600
rect 29698 15544 29703 15600
rect 12804 15542 29703 15544
rect 6361 15539 6427 15542
rect 7557 15539 7623 15542
rect 12525 15539 12591 15542
rect 29637 15539 29703 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 3417 15466 3483 15469
rect 11278 15466 11284 15468
rect 3417 15464 11284 15466
rect 3417 15408 3422 15464
rect 3478 15408 11284 15464
rect 3417 15406 11284 15408
rect 3417 15403 3483 15406
rect 11278 15404 11284 15406
rect 11348 15404 11354 15468
rect 12157 15466 12223 15469
rect 26233 15466 26299 15469
rect 12157 15464 26299 15466
rect 12157 15408 12162 15464
rect 12218 15408 26238 15464
rect 26294 15408 26299 15464
rect 12157 15406 26299 15408
rect 12157 15403 12223 15406
rect 26233 15403 26299 15406
rect 4337 15332 4403 15333
rect 13537 15332 13603 15333
rect 15009 15332 15075 15333
rect 4286 15268 4292 15332
rect 4356 15330 4403 15332
rect 13486 15330 13492 15332
rect 4356 15328 4448 15330
rect 4398 15272 4448 15328
rect 4356 15270 4448 15272
rect 13446 15270 13492 15330
rect 13556 15328 13603 15332
rect 14958 15330 14964 15332
rect 13598 15272 13603 15328
rect 4356 15268 4403 15270
rect 13486 15268 13492 15270
rect 13556 15268 13603 15272
rect 14918 15270 14964 15330
rect 15028 15328 15075 15332
rect 15070 15272 15075 15328
rect 14958 15268 14964 15270
rect 15028 15268 15075 15272
rect 4337 15267 4403 15268
rect 13537 15267 13603 15268
rect 15009 15267 15075 15268
rect 19149 15330 19215 15333
rect 23657 15330 23723 15333
rect 19149 15328 23723 15330
rect 19149 15272 19154 15328
rect 19210 15272 23662 15328
rect 23718 15272 23723 15328
rect 19149 15270 23723 15272
rect 19149 15267 19215 15270
rect 23657 15267 23723 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 9070 15132 9076 15196
rect 9140 15194 9146 15196
rect 10133 15194 10199 15197
rect 9140 15192 10199 15194
rect 9140 15136 10138 15192
rect 10194 15136 10199 15192
rect 9140 15134 10199 15136
rect 9140 15132 9146 15134
rect 10133 15131 10199 15134
rect 11973 15194 12039 15197
rect 13905 15194 13971 15197
rect 11973 15192 13971 15194
rect 11973 15136 11978 15192
rect 12034 15136 13910 15192
rect 13966 15136 13971 15192
rect 11973 15134 13971 15136
rect 11973 15131 12039 15134
rect 13905 15131 13971 15134
rect 14089 15194 14155 15197
rect 19977 15194 20043 15197
rect 25589 15194 25655 15197
rect 27613 15194 27679 15197
rect 14089 15192 14290 15194
rect 14089 15136 14094 15192
rect 14150 15136 14290 15192
rect 14089 15134 14290 15136
rect 14089 15131 14155 15134
rect 0 15058 800 15088
rect 1117 15058 1183 15061
rect 0 15056 1183 15058
rect 0 15000 1122 15056
rect 1178 15000 1183 15056
rect 0 14998 1183 15000
rect 0 14968 800 14998
rect 1117 14995 1183 14998
rect 5993 15058 6059 15061
rect 14230 15058 14290 15134
rect 19977 15192 27679 15194
rect 19977 15136 19982 15192
rect 20038 15136 25594 15192
rect 25650 15136 27618 15192
rect 27674 15136 27679 15192
rect 19977 15134 27679 15136
rect 19977 15131 20043 15134
rect 25589 15131 25655 15134
rect 27613 15131 27679 15134
rect 22553 15058 22619 15061
rect 5993 15056 14106 15058
rect 5993 15000 5998 15056
rect 6054 15000 14106 15056
rect 5993 14998 14106 15000
rect 14230 15056 22619 15058
rect 14230 15000 22558 15056
rect 22614 15000 22619 15056
rect 14230 14998 22619 15000
rect 5993 14995 6059 14998
rect 3734 14860 3740 14924
rect 3804 14922 3810 14924
rect 13905 14922 13971 14925
rect 3804 14920 13971 14922
rect 3804 14864 13910 14920
rect 13966 14864 13971 14920
rect 3804 14862 13971 14864
rect 14046 14922 14106 14998
rect 22553 14995 22619 14998
rect 21173 14922 21239 14925
rect 14046 14920 21239 14922
rect 14046 14864 21178 14920
rect 21234 14864 21239 14920
rect 14046 14862 21239 14864
rect 3804 14860 3810 14862
rect 13905 14859 13971 14862
rect 21173 14859 21239 14862
rect 5574 14724 5580 14788
rect 5644 14786 5650 14788
rect 10685 14786 10751 14789
rect 10961 14786 11027 14789
rect 5644 14784 11027 14786
rect 5644 14728 10690 14784
rect 10746 14728 10966 14784
rect 11022 14728 11027 14784
rect 5644 14726 11027 14728
rect 5644 14724 5650 14726
rect 10685 14723 10751 14726
rect 10961 14723 11027 14726
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 8477 14650 8543 14653
rect 8886 14650 8892 14652
rect 8477 14648 8892 14650
rect 8477 14592 8482 14648
rect 8538 14592 8892 14648
rect 8477 14590 8892 14592
rect 8477 14587 8543 14590
rect 8886 14588 8892 14590
rect 8956 14588 8962 14652
rect 9765 14650 9831 14653
rect 12801 14650 12867 14653
rect 9765 14648 12867 14650
rect 9765 14592 9770 14648
rect 9826 14592 12806 14648
rect 12862 14592 12867 14648
rect 9765 14590 12867 14592
rect 9765 14587 9831 14590
rect 12801 14587 12867 14590
rect 3601 14514 3667 14517
rect 11697 14514 11763 14517
rect 3601 14512 11763 14514
rect 3601 14456 3606 14512
rect 3662 14456 11702 14512
rect 11758 14456 11763 14512
rect 3601 14454 11763 14456
rect 3601 14451 3667 14454
rect 11697 14451 11763 14454
rect 11973 14514 12039 14517
rect 12249 14514 12315 14517
rect 11973 14512 12315 14514
rect 11973 14456 11978 14512
rect 12034 14456 12254 14512
rect 12310 14456 12315 14512
rect 11973 14454 12315 14456
rect 11973 14451 12039 14454
rect 12249 14451 12315 14454
rect 16849 14514 16915 14517
rect 24945 14514 25011 14517
rect 16849 14512 25011 14514
rect 16849 14456 16854 14512
rect 16910 14456 24950 14512
rect 25006 14456 25011 14512
rect 16849 14454 25011 14456
rect 16849 14451 16915 14454
rect 24945 14451 25011 14454
rect 7598 14316 7604 14380
rect 7668 14378 7674 14380
rect 8201 14378 8267 14381
rect 7668 14376 8267 14378
rect 7668 14320 8206 14376
rect 8262 14320 8267 14376
rect 7668 14318 8267 14320
rect 7668 14316 7674 14318
rect 8201 14315 8267 14318
rect 8845 14380 8911 14381
rect 8845 14376 8892 14380
rect 8956 14378 8962 14380
rect 10133 14378 10199 14381
rect 12709 14378 12775 14381
rect 8845 14320 8850 14376
rect 8845 14316 8892 14320
rect 8956 14318 9002 14378
rect 10133 14376 12775 14378
rect 10133 14320 10138 14376
rect 10194 14320 12714 14376
rect 12770 14320 12775 14376
rect 10133 14318 12775 14320
rect 8956 14316 8962 14318
rect 8845 14315 8911 14316
rect 10133 14315 10199 14318
rect 12709 14315 12775 14318
rect 15193 14378 15259 14381
rect 20069 14378 20135 14381
rect 15193 14376 20135 14378
rect 15193 14320 15198 14376
rect 15254 14320 20074 14376
rect 20130 14320 20135 14376
rect 15193 14318 20135 14320
rect 15193 14315 15259 14318
rect 20069 14315 20135 14318
rect 20345 14378 20411 14381
rect 34697 14378 34763 14381
rect 20345 14376 34763 14378
rect 20345 14320 20350 14376
rect 20406 14320 34702 14376
rect 34758 14320 34763 14376
rect 20345 14318 34763 14320
rect 20345 14315 20411 14318
rect 34697 14315 34763 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 8334 14180 8340 14244
rect 8404 14242 8410 14244
rect 13905 14242 13971 14245
rect 8404 14240 13971 14242
rect 8404 14184 13910 14240
rect 13966 14184 13971 14240
rect 8404 14182 13971 14184
rect 8404 14180 8410 14182
rect 13905 14179 13971 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 11421 14106 11487 14109
rect 13353 14106 13419 14109
rect 11421 14104 13419 14106
rect 11421 14048 11426 14104
rect 11482 14048 13358 14104
rect 13414 14048 13419 14104
rect 11421 14046 13419 14048
rect 11421 14043 11487 14046
rect 13353 14043 13419 14046
rect 15653 14106 15719 14109
rect 17217 14106 17283 14109
rect 15653 14104 17283 14106
rect 15653 14048 15658 14104
rect 15714 14048 17222 14104
rect 17278 14048 17283 14104
rect 15653 14046 17283 14048
rect 15653 14043 15719 14046
rect 17217 14043 17283 14046
rect 20253 14106 20319 14109
rect 24117 14106 24183 14109
rect 20253 14104 24183 14106
rect 20253 14048 20258 14104
rect 20314 14048 24122 14104
rect 24178 14048 24183 14104
rect 20253 14046 24183 14048
rect 20253 14043 20319 14046
rect 24117 14043 24183 14046
rect 3509 13970 3575 13973
rect 4429 13970 4495 13973
rect 11605 13970 11671 13973
rect 3509 13968 11671 13970
rect 3509 13912 3514 13968
rect 3570 13912 4434 13968
rect 4490 13912 11610 13968
rect 11666 13912 11671 13968
rect 3509 13910 11671 13912
rect 3509 13907 3575 13910
rect 4429 13907 4495 13910
rect 11605 13907 11671 13910
rect 12157 13970 12223 13973
rect 33685 13970 33751 13973
rect 12157 13968 33751 13970
rect 12157 13912 12162 13968
rect 12218 13912 33690 13968
rect 33746 13912 33751 13968
rect 12157 13910 33751 13912
rect 12157 13907 12223 13910
rect 33685 13907 33751 13910
rect 0 13834 800 13864
rect 2037 13834 2103 13837
rect 5533 13836 5599 13837
rect 5533 13834 5580 13836
rect 0 13832 2103 13834
rect 0 13776 2042 13832
rect 2098 13776 2103 13832
rect 0 13774 2103 13776
rect 5488 13832 5580 13834
rect 5488 13776 5538 13832
rect 5488 13774 5580 13776
rect 0 13744 800 13774
rect 2037 13771 2103 13774
rect 5533 13772 5580 13774
rect 5644 13772 5650 13836
rect 9581 13834 9647 13837
rect 10961 13834 11027 13837
rect 9581 13832 11027 13834
rect 9581 13776 9586 13832
rect 9642 13776 10966 13832
rect 11022 13776 11027 13832
rect 9581 13774 11027 13776
rect 5533 13771 5599 13772
rect 9581 13771 9647 13774
rect 10961 13771 11027 13774
rect 12893 13834 12959 13837
rect 32857 13834 32923 13837
rect 12893 13832 32923 13834
rect 12893 13776 12898 13832
rect 12954 13776 32862 13832
rect 32918 13776 32923 13832
rect 12893 13774 32923 13776
rect 12893 13771 12959 13774
rect 32857 13771 32923 13774
rect 4889 13698 4955 13701
rect 5257 13700 5323 13701
rect 5022 13698 5028 13700
rect 4889 13696 5028 13698
rect 4889 13640 4894 13696
rect 4950 13640 5028 13696
rect 4889 13638 5028 13640
rect 4889 13635 4955 13638
rect 5022 13636 5028 13638
rect 5092 13636 5098 13700
rect 5206 13698 5212 13700
rect 5166 13638 5212 13698
rect 5276 13696 5323 13700
rect 5318 13640 5323 13696
rect 5206 13636 5212 13638
rect 5276 13636 5323 13640
rect 5257 13635 5323 13636
rect 10041 13698 10107 13701
rect 12198 13698 12204 13700
rect 10041 13696 12204 13698
rect 10041 13640 10046 13696
rect 10102 13640 12204 13696
rect 10041 13638 12204 13640
rect 10041 13635 10107 13638
rect 12198 13636 12204 13638
rect 12268 13636 12274 13700
rect 12801 13698 12867 13701
rect 12390 13696 12867 13698
rect 12390 13640 12806 13696
rect 12862 13640 12867 13696
rect 12390 13638 12867 13640
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 3366 13500 3372 13564
rect 3436 13562 3442 13564
rect 3601 13562 3667 13565
rect 12390 13562 12450 13638
rect 12801 13635 12867 13638
rect 26877 13698 26943 13701
rect 31753 13698 31819 13701
rect 26877 13696 31819 13698
rect 26877 13640 26882 13696
rect 26938 13640 31758 13696
rect 31814 13640 31819 13696
rect 26877 13638 31819 13640
rect 26877 13635 26943 13638
rect 31753 13635 31819 13638
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 3436 13560 12450 13562
rect 3436 13504 3606 13560
rect 3662 13504 12450 13560
rect 3436 13502 12450 13504
rect 13353 13562 13419 13565
rect 18045 13562 18111 13565
rect 18413 13562 18479 13565
rect 13353 13560 17050 13562
rect 13353 13504 13358 13560
rect 13414 13504 17050 13560
rect 13353 13502 17050 13504
rect 3436 13500 3442 13502
rect 3601 13499 3667 13502
rect 13353 13499 13419 13502
rect 0 13426 800 13456
rect 1117 13426 1183 13429
rect 0 13424 1183 13426
rect 0 13368 1122 13424
rect 1178 13368 1183 13424
rect 0 13366 1183 13368
rect 0 13336 800 13366
rect 1117 13363 1183 13366
rect 1761 13426 1827 13429
rect 1894 13426 1900 13428
rect 1761 13424 1900 13426
rect 1761 13368 1766 13424
rect 1822 13368 1900 13424
rect 1761 13366 1900 13368
rect 1761 13363 1827 13366
rect 1894 13364 1900 13366
rect 1964 13426 1970 13428
rect 14774 13426 14780 13428
rect 1964 13366 14780 13426
rect 1964 13364 1970 13366
rect 14774 13364 14780 13366
rect 14844 13364 14850 13428
rect 16990 13426 17050 13502
rect 18045 13560 18479 13562
rect 18045 13504 18050 13560
rect 18106 13504 18418 13560
rect 18474 13504 18479 13560
rect 18045 13502 18479 13504
rect 18045 13499 18111 13502
rect 18413 13499 18479 13502
rect 18781 13562 18847 13565
rect 22277 13562 22343 13565
rect 18781 13560 22343 13562
rect 18781 13504 18786 13560
rect 18842 13504 22282 13560
rect 22338 13504 22343 13560
rect 18781 13502 22343 13504
rect 18781 13499 18847 13502
rect 22277 13499 22343 13502
rect 23381 13562 23447 13565
rect 23749 13562 23815 13565
rect 23381 13560 23815 13562
rect 23381 13504 23386 13560
rect 23442 13504 23754 13560
rect 23810 13504 23815 13560
rect 23381 13502 23815 13504
rect 23381 13499 23447 13502
rect 23749 13499 23815 13502
rect 18638 13426 18644 13428
rect 16990 13366 18644 13426
rect 18638 13364 18644 13366
rect 18708 13364 18714 13428
rect 19742 13364 19748 13428
rect 19812 13426 19818 13428
rect 37641 13426 37707 13429
rect 19812 13424 37707 13426
rect 19812 13368 37646 13424
rect 37702 13368 37707 13424
rect 19812 13366 37707 13368
rect 19812 13364 19818 13366
rect 37641 13363 37707 13366
rect 4429 13290 4495 13293
rect 4429 13288 9690 13290
rect 4429 13232 4434 13288
rect 4490 13232 9690 13288
rect 4429 13230 9690 13232
rect 4429 13227 4495 13230
rect 4981 13154 5047 13157
rect 7189 13154 7255 13157
rect 4981 13152 7255 13154
rect 4981 13096 4986 13152
rect 5042 13096 7194 13152
rect 7250 13096 7255 13152
rect 4981 13094 7255 13096
rect 9630 13154 9690 13230
rect 10910 13228 10916 13292
rect 10980 13290 10986 13292
rect 37089 13290 37155 13293
rect 10980 13288 37155 13290
rect 10980 13232 37094 13288
rect 37150 13232 37155 13288
rect 10980 13230 37155 13232
rect 10980 13228 10986 13230
rect 37089 13227 37155 13230
rect 9990 13154 9996 13156
rect 9630 13094 9996 13154
rect 4981 13091 5047 13094
rect 7189 13091 7255 13094
rect 9990 13092 9996 13094
rect 10060 13154 10066 13156
rect 14089 13154 14155 13157
rect 10060 13152 14155 13154
rect 10060 13096 14094 13152
rect 14150 13096 14155 13152
rect 10060 13094 14155 13096
rect 10060 13092 10066 13094
rect 14089 13091 14155 13094
rect 19926 13092 19932 13156
rect 19996 13154 20002 13156
rect 26877 13154 26943 13157
rect 19996 13152 26943 13154
rect 19996 13096 26882 13152
rect 26938 13096 26943 13152
rect 19996 13094 26943 13096
rect 19996 13092 20002 13094
rect 26877 13091 26943 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 3233 13018 3299 13021
rect 0 13016 3299 13018
rect 0 12960 3238 13016
rect 3294 12960 3299 13016
rect 0 12958 3299 12960
rect 0 12928 800 12958
rect 3233 12955 3299 12958
rect 9254 12956 9260 13020
rect 9324 13018 9330 13020
rect 10225 13018 10291 13021
rect 12709 13020 12775 13021
rect 12709 13018 12756 13020
rect 9324 13016 10291 13018
rect 9324 12960 10230 13016
rect 10286 12960 10291 13016
rect 9324 12958 10291 12960
rect 12664 13016 12756 13018
rect 12820 13018 12826 13020
rect 13353 13018 13419 13021
rect 12820 13016 13419 13018
rect 12664 12960 12714 13016
rect 12820 12960 13358 13016
rect 13414 12960 13419 13016
rect 12664 12958 12756 12960
rect 9324 12956 9330 12958
rect 10225 12955 10291 12958
rect 12709 12956 12756 12958
rect 12820 12958 13419 12960
rect 12820 12956 12826 12958
rect 12709 12955 12775 12956
rect 13353 12955 13419 12958
rect 13537 13018 13603 13021
rect 13670 13018 13676 13020
rect 13537 13016 13676 13018
rect 13537 12960 13542 13016
rect 13598 12960 13676 13016
rect 13537 12958 13676 12960
rect 13537 12955 13603 12958
rect 13670 12956 13676 12958
rect 13740 12956 13746 13020
rect 4061 12882 4127 12885
rect 5349 12882 5415 12885
rect 4061 12880 5415 12882
rect 4061 12824 4066 12880
rect 4122 12824 5354 12880
rect 5410 12824 5415 12880
rect 4061 12822 5415 12824
rect 4061 12819 4127 12822
rect 5349 12819 5415 12822
rect 5942 12820 5948 12884
rect 6012 12882 6018 12884
rect 6085 12882 6151 12885
rect 6012 12880 6151 12882
rect 6012 12824 6090 12880
rect 6146 12824 6151 12880
rect 6012 12822 6151 12824
rect 6012 12820 6018 12822
rect 6085 12819 6151 12822
rect 6269 12882 6335 12885
rect 11973 12882 12039 12885
rect 6269 12880 12039 12882
rect 6269 12824 6274 12880
rect 6330 12824 11978 12880
rect 12034 12824 12039 12880
rect 6269 12822 12039 12824
rect 6269 12819 6335 12822
rect 11973 12819 12039 12822
rect 12985 12882 13051 12885
rect 19558 12882 19564 12884
rect 12985 12880 19564 12882
rect 12985 12824 12990 12880
rect 13046 12824 19564 12880
rect 12985 12822 19564 12824
rect 12985 12819 13051 12822
rect 19558 12820 19564 12822
rect 19628 12820 19634 12884
rect 19885 12882 19951 12885
rect 41505 12882 41571 12885
rect 19885 12880 41571 12882
rect 19885 12824 19890 12880
rect 19946 12824 41510 12880
rect 41566 12824 41571 12880
rect 19885 12822 41571 12824
rect 19885 12819 19951 12822
rect 41505 12819 41571 12822
rect 4613 12746 4679 12749
rect 2730 12744 4679 12746
rect 2730 12688 4618 12744
rect 4674 12688 4679 12744
rect 2730 12686 4679 12688
rect 0 12610 800 12640
rect 2730 12610 2790 12686
rect 4613 12683 4679 12686
rect 9990 12684 9996 12748
rect 10060 12746 10066 12748
rect 24209 12746 24275 12749
rect 10060 12744 24275 12746
rect 10060 12688 24214 12744
rect 24270 12688 24275 12744
rect 10060 12686 24275 12688
rect 10060 12684 10066 12686
rect 24209 12683 24275 12686
rect 0 12550 2790 12610
rect 3325 12610 3391 12613
rect 3601 12610 3667 12613
rect 11789 12610 11855 12613
rect 3325 12608 3434 12610
rect 3325 12552 3330 12608
rect 3386 12552 3434 12608
rect 0 12520 800 12550
rect 3325 12547 3434 12552
rect 3601 12608 11855 12610
rect 3601 12552 3606 12608
rect 3662 12552 11794 12608
rect 11850 12552 11855 12608
rect 3601 12550 11855 12552
rect 3601 12547 3667 12550
rect 11789 12547 11855 12550
rect 14181 12610 14247 12613
rect 14549 12610 14615 12613
rect 14181 12608 14615 12610
rect 14181 12552 14186 12608
rect 14242 12552 14554 12608
rect 14610 12552 14615 12608
rect 14181 12550 14615 12552
rect 14181 12547 14247 12550
rect 14549 12547 14615 12550
rect 14825 12610 14891 12613
rect 18689 12610 18755 12613
rect 14825 12608 18755 12610
rect 14825 12552 14830 12608
rect 14886 12552 18694 12608
rect 18750 12552 18755 12608
rect 14825 12550 18755 12552
rect 14825 12547 14891 12550
rect 18689 12547 18755 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 3374 12474 3434 12547
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 4061 12474 4127 12477
rect 3374 12472 4127 12474
rect 3374 12416 4066 12472
rect 4122 12416 4127 12472
rect 3374 12414 4127 12416
rect 4061 12411 4127 12414
rect 2497 12338 2563 12341
rect 4061 12338 4127 12341
rect 4337 12340 4403 12341
rect 4286 12338 4292 12340
rect 2497 12336 4127 12338
rect 2497 12280 2502 12336
rect 2558 12280 4066 12336
rect 4122 12280 4127 12336
rect 2497 12278 4127 12280
rect 4246 12278 4292 12338
rect 4356 12336 4403 12340
rect 4398 12280 4403 12336
rect 2497 12275 2563 12278
rect 4061 12275 4127 12278
rect 4286 12276 4292 12278
rect 4356 12276 4403 12280
rect 4337 12275 4403 12276
rect 5625 12338 5691 12341
rect 6361 12338 6427 12341
rect 5625 12336 6427 12338
rect 5625 12280 5630 12336
rect 5686 12280 6366 12336
rect 6422 12280 6427 12336
rect 5625 12278 6427 12280
rect 5625 12275 5691 12278
rect 6361 12275 6427 12278
rect 14641 12338 14707 12341
rect 35985 12338 36051 12341
rect 14641 12336 36051 12338
rect 14641 12280 14646 12336
rect 14702 12280 35990 12336
rect 36046 12280 36051 12336
rect 14641 12278 36051 12280
rect 14641 12275 14707 12278
rect 35985 12275 36051 12278
rect 0 12202 800 12232
rect 1761 12202 1827 12205
rect 0 12200 1827 12202
rect 0 12144 1766 12200
rect 1822 12144 1827 12200
rect 0 12142 1827 12144
rect 0 12112 800 12142
rect 1761 12139 1827 12142
rect 3233 12202 3299 12205
rect 8702 12202 8708 12204
rect 3233 12200 8708 12202
rect 3233 12144 3238 12200
rect 3294 12144 8708 12200
rect 3233 12142 8708 12144
rect 3233 12139 3299 12142
rect 8702 12140 8708 12142
rect 8772 12140 8778 12204
rect 11789 12202 11855 12205
rect 29545 12202 29611 12205
rect 11789 12200 29611 12202
rect 11789 12144 11794 12200
rect 11850 12144 29550 12200
rect 29606 12144 29611 12200
rect 11789 12142 29611 12144
rect 11789 12139 11855 12142
rect 29545 12139 29611 12142
rect 4286 12004 4292 12068
rect 4356 12066 4362 12068
rect 4429 12066 4495 12069
rect 4356 12064 4495 12066
rect 4356 12008 4434 12064
rect 4490 12008 4495 12064
rect 4356 12006 4495 12008
rect 4356 12004 4362 12006
rect 4429 12003 4495 12006
rect 4889 12066 4955 12069
rect 5349 12066 5415 12069
rect 6545 12066 6611 12069
rect 7373 12066 7439 12069
rect 4889 12064 7439 12066
rect 4889 12008 4894 12064
rect 4950 12008 5354 12064
rect 5410 12008 6550 12064
rect 6606 12008 7378 12064
rect 7434 12008 7439 12064
rect 4889 12006 7439 12008
rect 4889 12003 4955 12006
rect 5349 12003 5415 12006
rect 6545 12003 6611 12006
rect 7373 12003 7439 12006
rect 13997 12066 14063 12069
rect 15377 12066 15443 12069
rect 16297 12068 16363 12069
rect 16246 12066 16252 12068
rect 13997 12064 15443 12066
rect 13997 12008 14002 12064
rect 14058 12008 15382 12064
rect 15438 12008 15443 12064
rect 13997 12006 15443 12008
rect 16206 12006 16252 12066
rect 16316 12064 16363 12068
rect 16358 12008 16363 12064
rect 13997 12003 14063 12006
rect 15377 12003 15443 12006
rect 16246 12004 16252 12006
rect 16316 12004 16363 12008
rect 16297 12003 16363 12004
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 2405 11932 2471 11933
rect 2405 11930 2452 11932
rect 2360 11928 2452 11930
rect 2360 11872 2410 11928
rect 2360 11870 2452 11872
rect 2405 11868 2452 11870
rect 2516 11868 2522 11932
rect 11973 11930 12039 11933
rect 17493 11930 17559 11933
rect 11973 11928 17559 11930
rect 11973 11872 11978 11928
rect 12034 11872 17498 11928
rect 17554 11872 17559 11928
rect 11973 11870 17559 11872
rect 2405 11867 2471 11868
rect 11973 11867 12039 11870
rect 17493 11867 17559 11870
rect 0 11794 800 11824
rect 3734 11794 3740 11796
rect 0 11734 3740 11794
rect 0 11704 800 11734
rect 3734 11732 3740 11734
rect 3804 11732 3810 11796
rect 5390 11732 5396 11796
rect 5460 11794 5466 11796
rect 10501 11794 10567 11797
rect 5460 11792 10567 11794
rect 5460 11736 10506 11792
rect 10562 11736 10567 11792
rect 5460 11734 10567 11736
rect 5460 11732 5466 11734
rect 10501 11731 10567 11734
rect 11697 11794 11763 11797
rect 20805 11794 20871 11797
rect 25497 11794 25563 11797
rect 11697 11792 25563 11794
rect 11697 11736 11702 11792
rect 11758 11736 20810 11792
rect 20866 11736 25502 11792
rect 25558 11736 25563 11792
rect 11697 11734 25563 11736
rect 11697 11731 11763 11734
rect 20805 11731 20871 11734
rect 25497 11731 25563 11734
rect 1853 11658 1919 11661
rect 13169 11658 13235 11661
rect 1853 11656 13235 11658
rect 1853 11600 1858 11656
rect 1914 11600 13174 11656
rect 13230 11600 13235 11656
rect 1853 11598 13235 11600
rect 1853 11595 1919 11598
rect 13169 11595 13235 11598
rect 16941 11658 17007 11661
rect 30005 11658 30071 11661
rect 16941 11656 30071 11658
rect 16941 11600 16946 11656
rect 17002 11600 30010 11656
rect 30066 11600 30071 11656
rect 16941 11598 30071 11600
rect 16941 11595 17007 11598
rect 30005 11595 30071 11598
rect 9765 11522 9831 11525
rect 12065 11522 12131 11525
rect 9765 11520 12131 11522
rect 9765 11464 9770 11520
rect 9826 11464 12070 11520
rect 12126 11464 12131 11520
rect 9765 11462 12131 11464
rect 9765 11459 9831 11462
rect 12065 11459 12131 11462
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 3601 11386 3667 11389
rect 4654 11386 4660 11388
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 2730 11250 2790 11326
rect 3601 11384 4660 11386
rect 3601 11328 3606 11384
rect 3662 11328 4660 11384
rect 3601 11326 4660 11328
rect 3601 11323 3667 11326
rect 4654 11324 4660 11326
rect 4724 11324 4730 11388
rect 8109 11386 8175 11389
rect 12709 11386 12775 11389
rect 8109 11384 12775 11386
rect 8109 11328 8114 11384
rect 8170 11328 12714 11384
rect 12770 11328 12775 11384
rect 8109 11326 12775 11328
rect 8109 11323 8175 11326
rect 12709 11323 12775 11326
rect 13537 11386 13603 11389
rect 14181 11388 14247 11389
rect 13670 11386 13676 11388
rect 13537 11384 13676 11386
rect 13537 11328 13542 11384
rect 13598 11328 13676 11384
rect 13537 11326 13676 11328
rect 13537 11323 13603 11326
rect 13670 11324 13676 11326
rect 13740 11324 13746 11388
rect 14181 11386 14228 11388
rect 14136 11384 14228 11386
rect 14136 11328 14186 11384
rect 14136 11326 14228 11328
rect 14181 11324 14228 11326
rect 14292 11324 14298 11388
rect 14181 11323 14247 11324
rect 3693 11250 3759 11253
rect 2730 11248 3759 11250
rect 2730 11192 3698 11248
rect 3754 11192 3759 11248
rect 2730 11190 3759 11192
rect 3693 11187 3759 11190
rect 7281 11250 7347 11253
rect 10501 11250 10567 11253
rect 18454 11250 18460 11252
rect 7281 11248 10242 11250
rect 7281 11192 7286 11248
rect 7342 11192 10242 11248
rect 7281 11190 10242 11192
rect 7281 11187 7347 11190
rect 1577 11114 1643 11117
rect 2037 11114 2103 11117
rect 9990 11114 9996 11116
rect 1577 11112 9996 11114
rect 1577 11056 1582 11112
rect 1638 11056 2042 11112
rect 2098 11056 9996 11112
rect 1577 11054 9996 11056
rect 1577 11051 1643 11054
rect 2037 11051 2103 11054
rect 9990 11052 9996 11054
rect 10060 11052 10066 11116
rect 10182 11114 10242 11190
rect 10501 11248 18460 11250
rect 10501 11192 10506 11248
rect 10562 11192 18460 11248
rect 10501 11190 18460 11192
rect 10501 11187 10567 11190
rect 18454 11188 18460 11190
rect 18524 11188 18530 11252
rect 22461 11114 22527 11117
rect 10182 11112 22527 11114
rect 10182 11056 22466 11112
rect 22522 11056 22527 11112
rect 10182 11054 22527 11056
rect 22461 11051 22527 11054
rect 0 10978 800 11008
rect 1853 10980 1919 10981
rect 1853 10978 1900 10980
rect 0 10888 858 10978
rect 1808 10976 1900 10978
rect 1808 10920 1858 10976
rect 1808 10918 1900 10920
rect 1853 10916 1900 10918
rect 1964 10916 1970 10980
rect 5533 10978 5599 10981
rect 9765 10980 9831 10981
rect 7230 10978 7236 10980
rect 5533 10976 7236 10978
rect 5533 10920 5538 10976
rect 5594 10920 7236 10976
rect 5533 10918 7236 10920
rect 1853 10915 1919 10916
rect 5533 10915 5599 10918
rect 7230 10916 7236 10918
rect 7300 10916 7306 10980
rect 9765 10976 9812 10980
rect 9876 10978 9882 10980
rect 9765 10920 9770 10976
rect 9765 10916 9812 10920
rect 9876 10918 9922 10978
rect 9876 10916 9882 10918
rect 12566 10916 12572 10980
rect 12636 10978 12642 10980
rect 13629 10978 13695 10981
rect 12636 10976 13695 10978
rect 12636 10920 13634 10976
rect 13690 10920 13695 10976
rect 12636 10918 13695 10920
rect 12636 10916 12642 10918
rect 9765 10915 9831 10916
rect 13629 10915 13695 10918
rect 798 10842 858 10888
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 2865 10842 2931 10845
rect 798 10840 2931 10842
rect 798 10784 2870 10840
rect 2926 10784 2931 10840
rect 798 10782 2931 10784
rect 2865 10779 2931 10782
rect 3785 10842 3851 10845
rect 3918 10842 3924 10844
rect 3785 10840 3924 10842
rect 3785 10784 3790 10840
rect 3846 10784 3924 10840
rect 3785 10782 3924 10784
rect 3785 10779 3851 10782
rect 3918 10780 3924 10782
rect 3988 10780 3994 10844
rect 11145 10842 11211 10845
rect 13905 10842 13971 10845
rect 11145 10840 13971 10842
rect 11145 10784 11150 10840
rect 11206 10784 13910 10840
rect 13966 10784 13971 10840
rect 11145 10782 13971 10784
rect 11145 10779 11211 10782
rect 13905 10779 13971 10782
rect 933 10706 999 10709
rect 1342 10706 1348 10708
rect 933 10704 1348 10706
rect 933 10648 938 10704
rect 994 10648 1348 10704
rect 933 10646 1348 10648
rect 933 10643 999 10646
rect 1342 10644 1348 10646
rect 1412 10644 1418 10708
rect 1853 10706 1919 10709
rect 5942 10706 5948 10708
rect 1853 10704 5948 10706
rect 1853 10648 1858 10704
rect 1914 10648 5948 10704
rect 1853 10646 5948 10648
rect 1853 10643 1919 10646
rect 5942 10644 5948 10646
rect 6012 10644 6018 10708
rect 10593 10706 10659 10709
rect 11830 10706 11836 10708
rect 10593 10704 11836 10706
rect 10593 10648 10598 10704
rect 10654 10648 11836 10704
rect 10593 10646 11836 10648
rect 10593 10643 10659 10646
rect 11830 10644 11836 10646
rect 11900 10644 11906 10708
rect 0 10570 800 10600
rect 3417 10570 3483 10573
rect 0 10568 3483 10570
rect 0 10512 3422 10568
rect 3478 10512 3483 10568
rect 0 10510 3483 10512
rect 0 10480 800 10510
rect 3417 10507 3483 10510
rect 15929 10570 15995 10573
rect 21909 10570 21975 10573
rect 15929 10568 21975 10570
rect 15929 10512 15934 10568
rect 15990 10512 21914 10568
rect 21970 10512 21975 10568
rect 15929 10510 21975 10512
rect 15929 10507 15995 10510
rect 21909 10507 21975 10510
rect 2405 10434 2471 10437
rect 2630 10434 2636 10436
rect 2405 10432 2636 10434
rect 2405 10376 2410 10432
rect 2466 10376 2636 10432
rect 2405 10374 2636 10376
rect 2405 10371 2471 10374
rect 2630 10372 2636 10374
rect 2700 10372 2706 10436
rect 7373 10434 7439 10437
rect 9254 10434 9260 10436
rect 7373 10432 9260 10434
rect 7373 10376 7378 10432
rect 7434 10376 9260 10432
rect 7373 10374 9260 10376
rect 7373 10371 7439 10374
rect 9254 10372 9260 10374
rect 9324 10372 9330 10436
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 3601 10162 3667 10165
rect 0 10160 3667 10162
rect 0 10104 3606 10160
rect 3662 10104 3667 10160
rect 0 10102 3667 10104
rect 0 10072 800 10102
rect 3601 10099 3667 10102
rect 4705 10162 4771 10165
rect 15326 10162 15332 10164
rect 4705 10160 15332 10162
rect 4705 10104 4710 10160
rect 4766 10104 15332 10160
rect 4705 10102 15332 10104
rect 4705 10099 4771 10102
rect 15326 10100 15332 10102
rect 15396 10100 15402 10164
rect 2957 10026 3023 10029
rect 3550 10026 3556 10028
rect 2957 10024 3556 10026
rect 2957 9968 2962 10024
rect 3018 9968 3556 10024
rect 2957 9966 3556 9968
rect 2957 9963 3023 9966
rect 3550 9964 3556 9966
rect 3620 10026 3626 10028
rect 35065 10026 35131 10029
rect 3620 10024 35131 10026
rect 3620 9968 35070 10024
rect 35126 9968 35131 10024
rect 3620 9966 35131 9968
rect 3620 9964 3626 9966
rect 35065 9963 35131 9966
rect 4521 9892 4587 9893
rect 4470 9890 4476 9892
rect 4430 9830 4476 9890
rect 4540 9888 4587 9892
rect 10501 9890 10567 9893
rect 4582 9832 4587 9888
rect 4470 9828 4476 9830
rect 4540 9828 4587 9832
rect 4521 9827 4587 9828
rect 8342 9888 10567 9890
rect 8342 9832 10506 9888
rect 10562 9832 10567 9888
rect 8342 9830 10567 9832
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 3509 9754 3575 9757
rect 5809 9756 5875 9757
rect 0 9752 3575 9754
rect 0 9696 3514 9752
rect 3570 9696 3575 9752
rect 0 9694 3575 9696
rect 0 9664 800 9694
rect 3509 9691 3575 9694
rect 5758 9692 5764 9756
rect 5828 9754 5875 9756
rect 5993 9754 6059 9757
rect 6126 9754 6132 9756
rect 5828 9752 5920 9754
rect 5870 9696 5920 9752
rect 5828 9694 5920 9696
rect 5993 9752 6132 9754
rect 5993 9696 5998 9752
rect 6054 9696 6132 9752
rect 5993 9694 6132 9696
rect 5828 9692 5875 9694
rect 5809 9691 5875 9692
rect 5993 9691 6059 9694
rect 6126 9692 6132 9694
rect 6196 9692 6202 9756
rect 6269 9754 6335 9757
rect 6678 9754 6684 9756
rect 6269 9752 6684 9754
rect 6269 9696 6274 9752
rect 6330 9696 6684 9752
rect 6269 9694 6684 9696
rect 6269 9691 6335 9694
rect 6678 9692 6684 9694
rect 6748 9692 6754 9756
rect 1485 9620 1551 9621
rect 3325 9620 3391 9621
rect 1485 9618 1532 9620
rect 1440 9616 1532 9618
rect 1440 9560 1490 9616
rect 1440 9558 1532 9560
rect 1485 9556 1532 9558
rect 1596 9556 1602 9620
rect 3325 9618 3372 9620
rect 3280 9616 3372 9618
rect 3280 9560 3330 9616
rect 3280 9558 3372 9560
rect 3325 9556 3372 9558
rect 3436 9556 3442 9620
rect 3969 9618 4035 9621
rect 4102 9618 4108 9620
rect 3969 9616 4108 9618
rect 3969 9560 3974 9616
rect 4030 9560 4108 9616
rect 3969 9558 4108 9560
rect 1485 9555 1551 9556
rect 3325 9555 3391 9556
rect 3969 9555 4035 9558
rect 4102 9556 4108 9558
rect 4172 9556 4178 9620
rect 7005 9618 7071 9621
rect 8342 9618 8402 9830
rect 10501 9827 10567 9830
rect 12157 9890 12223 9893
rect 13261 9890 13327 9893
rect 12157 9888 13327 9890
rect 12157 9832 12162 9888
rect 12218 9832 13266 9888
rect 13322 9832 13327 9888
rect 12157 9830 13327 9832
rect 12157 9827 12223 9830
rect 13261 9827 13327 9830
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 8937 9754 9003 9757
rect 9857 9754 9923 9757
rect 10685 9756 10751 9757
rect 10685 9754 10732 9756
rect 8937 9752 9923 9754
rect 8937 9696 8942 9752
rect 8998 9696 9862 9752
rect 9918 9696 9923 9752
rect 8937 9694 9923 9696
rect 10640 9752 10732 9754
rect 10640 9696 10690 9752
rect 10640 9694 10732 9696
rect 8937 9691 9003 9694
rect 9857 9691 9923 9694
rect 10685 9692 10732 9694
rect 10796 9692 10802 9756
rect 12750 9692 12756 9756
rect 12820 9754 12826 9756
rect 14958 9754 14964 9756
rect 12820 9694 14964 9754
rect 12820 9692 12826 9694
rect 14958 9692 14964 9694
rect 15028 9692 15034 9756
rect 10685 9691 10751 9692
rect 7005 9616 8402 9618
rect 7005 9560 7010 9616
rect 7066 9560 8402 9616
rect 7005 9558 8402 9560
rect 10317 9618 10383 9621
rect 13261 9618 13327 9621
rect 10317 9616 13327 9618
rect 10317 9560 10322 9616
rect 10378 9560 13266 9616
rect 13322 9560 13327 9616
rect 10317 9558 13327 9560
rect 7005 9555 7071 9558
rect 10317 9555 10383 9558
rect 13261 9555 13327 9558
rect 14038 9556 14044 9620
rect 14108 9618 14114 9620
rect 14181 9618 14247 9621
rect 14108 9616 14247 9618
rect 14108 9560 14186 9616
rect 14242 9560 14247 9616
rect 14108 9558 14247 9560
rect 14108 9556 14114 9558
rect 14181 9555 14247 9558
rect 15142 9556 15148 9620
rect 15212 9618 15218 9620
rect 36537 9618 36603 9621
rect 15212 9616 36603 9618
rect 15212 9560 36542 9616
rect 36598 9560 36603 9616
rect 15212 9558 36603 9560
rect 15212 9556 15218 9558
rect 36537 9555 36603 9558
rect 974 9420 980 9484
rect 1044 9482 1050 9484
rect 3417 9482 3483 9485
rect 1044 9480 3483 9482
rect 1044 9424 3422 9480
rect 3478 9424 3483 9480
rect 1044 9422 3483 9424
rect 1044 9420 1050 9422
rect 3417 9419 3483 9422
rect 4245 9482 4311 9485
rect 35157 9482 35223 9485
rect 4245 9480 35223 9482
rect 4245 9424 4250 9480
rect 4306 9424 35162 9480
rect 35218 9424 35223 9480
rect 4245 9422 35223 9424
rect 4245 9419 4311 9422
rect 35157 9419 35223 9422
rect 0 9346 800 9376
rect 2773 9346 2839 9349
rect 0 9344 2839 9346
rect 0 9288 2778 9344
rect 2834 9288 2839 9344
rect 0 9286 2839 9288
rect 0 9256 800 9286
rect 2773 9283 2839 9286
rect 6913 9346 6979 9349
rect 11421 9346 11487 9349
rect 6913 9344 11487 9346
rect 6913 9288 6918 9344
rect 6974 9288 11426 9344
rect 11482 9288 11487 9344
rect 6913 9286 11487 9288
rect 6913 9283 6979 9286
rect 11421 9283 11487 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 3877 9210 3943 9213
rect 12750 9210 12756 9212
rect 3877 9208 12756 9210
rect 3877 9152 3882 9208
rect 3938 9152 12756 9208
rect 3877 9150 12756 9152
rect 3877 9147 3943 9150
rect 12750 9148 12756 9150
rect 12820 9148 12826 9212
rect 3734 9012 3740 9076
rect 3804 9074 3810 9076
rect 3877 9074 3943 9077
rect 3804 9072 3943 9074
rect 3804 9016 3882 9072
rect 3938 9016 3943 9072
rect 3804 9014 3943 9016
rect 3804 9012 3810 9014
rect 3877 9011 3943 9014
rect 5165 9074 5231 9077
rect 5390 9074 5396 9076
rect 5165 9072 5396 9074
rect 5165 9016 5170 9072
rect 5226 9016 5396 9072
rect 5165 9014 5396 9016
rect 5165 9011 5231 9014
rect 5390 9012 5396 9014
rect 5460 9012 5466 9076
rect 5901 9074 5967 9077
rect 9438 9074 9444 9076
rect 5901 9072 9444 9074
rect 5901 9016 5906 9072
rect 5962 9016 9444 9072
rect 5901 9014 9444 9016
rect 5901 9011 5967 9014
rect 9438 9012 9444 9014
rect 9508 9012 9514 9076
rect 9673 9074 9739 9077
rect 10358 9074 10364 9076
rect 9673 9072 10364 9074
rect 9673 9016 9678 9072
rect 9734 9016 10364 9072
rect 9673 9014 10364 9016
rect 9673 9011 9739 9014
rect 10358 9012 10364 9014
rect 10428 9012 10434 9076
rect 10685 9074 10751 9077
rect 10961 9074 11027 9077
rect 10685 9072 11027 9074
rect 10685 9016 10690 9072
rect 10746 9016 10966 9072
rect 11022 9016 11027 9072
rect 10685 9014 11027 9016
rect 10685 9011 10751 9014
rect 10961 9011 11027 9014
rect 13169 9074 13235 9077
rect 24301 9074 24367 9077
rect 13169 9072 24367 9074
rect 13169 9016 13174 9072
rect 13230 9016 24306 9072
rect 24362 9016 24367 9072
rect 13169 9014 24367 9016
rect 13169 9011 13235 9014
rect 24301 9011 24367 9014
rect 0 8938 800 8968
rect 3141 8938 3207 8941
rect 0 8936 3207 8938
rect 0 8880 3146 8936
rect 3202 8880 3207 8936
rect 0 8878 3207 8880
rect 0 8848 800 8878
rect 3141 8875 3207 8878
rect 4245 8938 4311 8941
rect 36445 8938 36511 8941
rect 4245 8936 36511 8938
rect 4245 8880 4250 8936
rect 4306 8880 36450 8936
rect 36506 8880 36511 8936
rect 4245 8878 36511 8880
rect 4245 8875 4311 8878
rect 36445 8875 36511 8878
rect 10317 8802 10383 8805
rect 15142 8802 15148 8804
rect 10317 8800 15148 8802
rect 10317 8744 10322 8800
rect 10378 8744 15148 8800
rect 10317 8742 15148 8744
rect 10317 8739 10383 8742
rect 15142 8740 15148 8742
rect 15212 8740 15218 8804
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 11053 8668 11119 8669
rect 11053 8664 11100 8668
rect 11164 8666 11170 8668
rect 11329 8666 11395 8669
rect 11605 8668 11671 8669
rect 11462 8666 11468 8668
rect 11053 8608 11058 8664
rect 11053 8604 11100 8608
rect 11164 8606 11210 8666
rect 11329 8664 11468 8666
rect 11329 8608 11334 8664
rect 11390 8608 11468 8664
rect 11329 8606 11468 8608
rect 11164 8604 11170 8606
rect 11053 8603 11119 8604
rect 11329 8603 11395 8606
rect 11462 8604 11468 8606
rect 11532 8604 11538 8668
rect 11605 8664 11652 8668
rect 11716 8666 11722 8668
rect 12801 8666 12867 8669
rect 15469 8666 15535 8669
rect 11605 8608 11610 8664
rect 11605 8604 11652 8608
rect 11716 8606 11762 8666
rect 12801 8664 15535 8666
rect 12801 8608 12806 8664
rect 12862 8608 15474 8664
rect 15530 8608 15535 8664
rect 12801 8606 15535 8608
rect 11716 8604 11722 8606
rect 11605 8603 11671 8604
rect 12801 8603 12867 8606
rect 15469 8603 15535 8606
rect 0 8530 800 8560
rect 4797 8530 4863 8533
rect 0 8528 4863 8530
rect 0 8472 4802 8528
rect 4858 8472 4863 8528
rect 0 8470 4863 8472
rect 0 8440 800 8470
rect 4797 8467 4863 8470
rect 8293 8530 8359 8533
rect 9070 8530 9076 8532
rect 8293 8528 9076 8530
rect 8293 8472 8298 8528
rect 8354 8472 9076 8528
rect 8293 8470 9076 8472
rect 8293 8467 8359 8470
rect 9070 8468 9076 8470
rect 9140 8530 9146 8532
rect 9305 8530 9371 8533
rect 9140 8528 9371 8530
rect 9140 8472 9310 8528
rect 9366 8472 9371 8528
rect 9140 8470 9371 8472
rect 9140 8468 9146 8470
rect 9305 8467 9371 8470
rect 11145 8530 11211 8533
rect 15510 8530 15516 8532
rect 11145 8528 15516 8530
rect 11145 8472 11150 8528
rect 11206 8472 15516 8528
rect 11145 8470 15516 8472
rect 11145 8467 11211 8470
rect 15510 8468 15516 8470
rect 15580 8468 15586 8532
rect 8109 8394 8175 8397
rect 36721 8394 36787 8397
rect 8109 8392 36787 8394
rect 8109 8336 8114 8392
rect 8170 8336 36726 8392
rect 36782 8336 36787 8392
rect 8109 8334 36787 8336
rect 8109 8331 8175 8334
rect 36721 8331 36787 8334
rect 4889 8258 4955 8261
rect 5206 8258 5212 8260
rect 4889 8256 5212 8258
rect 4889 8200 4894 8256
rect 4950 8200 5212 8256
rect 4889 8198 5212 8200
rect 4889 8195 4955 8198
rect 5206 8196 5212 8198
rect 5276 8196 5282 8260
rect 6729 8258 6795 8261
rect 8477 8258 8543 8261
rect 6729 8256 8543 8258
rect 6729 8200 6734 8256
rect 6790 8200 8482 8256
rect 8538 8200 8543 8256
rect 6729 8198 8543 8200
rect 6729 8195 6795 8198
rect 8477 8195 8543 8198
rect 9857 8258 9923 8261
rect 12525 8258 12591 8261
rect 9857 8256 12591 8258
rect 9857 8200 9862 8256
rect 9918 8200 12530 8256
rect 12586 8200 12591 8256
rect 9857 8198 12591 8200
rect 9857 8195 9923 8198
rect 12525 8195 12591 8198
rect 13905 8258 13971 8261
rect 18505 8258 18571 8261
rect 13905 8256 18571 8258
rect 13905 8200 13910 8256
rect 13966 8200 18510 8256
rect 18566 8200 18571 8256
rect 13905 8198 18571 8200
rect 13905 8195 13971 8198
rect 18505 8195 18571 8198
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2313 8122 2379 8125
rect 0 8120 2379 8122
rect 0 8064 2318 8120
rect 2374 8064 2379 8120
rect 0 8062 2379 8064
rect 0 8032 800 8062
rect 2313 8059 2379 8062
rect 9857 8122 9923 8125
rect 10041 8122 10107 8125
rect 9857 8120 10107 8122
rect 9857 8064 9862 8120
rect 9918 8064 10046 8120
rect 10102 8064 10107 8120
rect 9857 8062 10107 8064
rect 9857 8059 9923 8062
rect 10041 8059 10107 8062
rect 12198 8060 12204 8124
rect 12268 8122 12274 8124
rect 12341 8122 12407 8125
rect 12268 8120 12407 8122
rect 12268 8064 12346 8120
rect 12402 8064 12407 8120
rect 12268 8062 12407 8064
rect 12268 8060 12274 8062
rect 12341 8059 12407 8062
rect 4705 7986 4771 7989
rect 9397 7986 9463 7989
rect 24761 7986 24827 7989
rect 4705 7984 8586 7986
rect 4705 7928 4710 7984
rect 4766 7928 8586 7984
rect 4705 7926 8586 7928
rect 4705 7923 4771 7926
rect 2773 7850 2839 7853
rect 8526 7850 8586 7926
rect 9397 7984 24827 7986
rect 9397 7928 9402 7984
rect 9458 7928 24766 7984
rect 24822 7928 24827 7984
rect 9397 7926 24827 7928
rect 9397 7923 9463 7926
rect 24761 7923 24827 7926
rect 22369 7850 22435 7853
rect 2773 7848 8402 7850
rect 2773 7792 2778 7848
rect 2834 7792 8402 7848
rect 2773 7790 8402 7792
rect 8526 7848 22435 7850
rect 8526 7792 22374 7848
rect 22430 7792 22435 7848
rect 8526 7790 22435 7792
rect 2773 7787 2839 7790
rect 0 7714 800 7744
rect 4337 7714 4403 7717
rect 0 7712 4403 7714
rect 0 7656 4342 7712
rect 4398 7656 4403 7712
rect 0 7654 4403 7656
rect 8342 7714 8402 7790
rect 22369 7787 22435 7790
rect 15694 7714 15700 7716
rect 8342 7654 15700 7714
rect 0 7624 800 7654
rect 4337 7651 4403 7654
rect 15694 7652 15700 7654
rect 15764 7652 15770 7716
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 1158 7516 1164 7580
rect 1228 7578 1234 7580
rect 4613 7578 4679 7581
rect 1228 7576 4679 7578
rect 1228 7520 4618 7576
rect 4674 7520 4679 7576
rect 1228 7518 4679 7520
rect 1228 7516 1234 7518
rect 4613 7515 4679 7518
rect 8661 7578 8727 7581
rect 8661 7576 17234 7578
rect 8661 7520 8666 7576
rect 8722 7520 17234 7576
rect 8661 7518 17234 7520
rect 8661 7515 8727 7518
rect 3233 7442 3299 7445
rect 7373 7444 7439 7445
rect 3550 7442 3556 7444
rect 3233 7440 3556 7442
rect 3233 7384 3238 7440
rect 3294 7384 3556 7440
rect 3233 7382 3556 7384
rect 3233 7379 3299 7382
rect 3550 7380 3556 7382
rect 3620 7380 3626 7444
rect 7373 7442 7420 7444
rect 7328 7440 7420 7442
rect 7328 7384 7378 7440
rect 7328 7382 7420 7384
rect 7373 7380 7420 7382
rect 7484 7380 7490 7444
rect 9857 7442 9923 7445
rect 11329 7442 11395 7445
rect 17174 7442 17234 7518
rect 36997 7442 37063 7445
rect 9857 7440 11395 7442
rect 9857 7384 9862 7440
rect 9918 7384 11334 7440
rect 11390 7384 11395 7440
rect 9857 7382 11395 7384
rect 7373 7379 7439 7380
rect 9857 7379 9923 7382
rect 11329 7379 11395 7382
rect 12574 7382 17050 7442
rect 17174 7440 37063 7442
rect 17174 7384 37002 7440
rect 37058 7384 37063 7440
rect 17174 7382 37063 7384
rect 0 7306 800 7336
rect 4521 7306 4587 7309
rect 0 7304 4587 7306
rect 0 7248 4526 7304
rect 4582 7248 4587 7304
rect 0 7246 4587 7248
rect 0 7216 800 7246
rect 4521 7243 4587 7246
rect 6821 7306 6887 7309
rect 12574 7306 12634 7382
rect 16990 7306 17050 7382
rect 36997 7379 37063 7382
rect 25129 7306 25195 7309
rect 6821 7304 12634 7306
rect 6821 7248 6826 7304
rect 6882 7248 12634 7304
rect 6821 7246 12634 7248
rect 12758 7246 16866 7306
rect 16990 7304 25195 7306
rect 16990 7248 25134 7304
rect 25190 7248 25195 7304
rect 16990 7246 25195 7248
rect 6821 7243 6887 7246
rect 6269 7170 6335 7173
rect 12758 7170 12818 7246
rect 6269 7168 12818 7170
rect 6269 7112 6274 7168
rect 6330 7112 12818 7168
rect 6269 7110 12818 7112
rect 13353 7170 13419 7173
rect 13670 7170 13676 7172
rect 13353 7168 13676 7170
rect 13353 7112 13358 7168
rect 13414 7112 13676 7168
rect 13353 7110 13676 7112
rect 6269 7107 6335 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 7192 7037 7252 7110
rect 13353 7107 13419 7110
rect 13670 7108 13676 7110
rect 13740 7108 13746 7172
rect 16806 7170 16866 7246
rect 25129 7243 25195 7246
rect 22737 7170 22803 7173
rect 16806 7168 22803 7170
rect 16806 7112 22742 7168
rect 22798 7112 22803 7168
rect 16806 7110 22803 7112
rect 22737 7107 22803 7110
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 7189 7032 7255 7037
rect 7189 6976 7194 7032
rect 7250 6976 7255 7032
rect 7189 6971 7255 6976
rect 9673 7034 9739 7037
rect 10174 7034 10180 7036
rect 9673 7032 10180 7034
rect 9673 6976 9678 7032
rect 9734 6976 10180 7032
rect 9673 6974 10180 6976
rect 9673 6971 9739 6974
rect 10174 6972 10180 6974
rect 10244 6972 10250 7036
rect 12341 7034 12407 7037
rect 22502 7034 22508 7036
rect 12341 7032 12818 7034
rect 12341 6976 12346 7032
rect 12402 6976 12818 7032
rect 12341 6974 12818 6976
rect 12341 6971 12407 6974
rect 0 6898 800 6928
rect 6913 6898 6979 6901
rect 8886 6898 8892 6900
rect 0 6838 2698 6898
rect 0 6808 800 6838
rect 2638 6762 2698 6838
rect 6913 6896 8892 6898
rect 6913 6840 6918 6896
rect 6974 6840 8892 6896
rect 6913 6838 8892 6840
rect 6913 6835 6979 6838
rect 8886 6836 8892 6838
rect 8956 6836 8962 6900
rect 12758 6898 12818 6974
rect 13494 6974 22508 7034
rect 13494 6898 13554 6974
rect 22502 6972 22508 6974
rect 22572 6972 22578 7036
rect 12758 6838 13554 6898
rect 3141 6762 3207 6765
rect 2638 6760 3207 6762
rect 2638 6704 3146 6760
rect 3202 6704 3207 6760
rect 2638 6702 3207 6704
rect 3141 6699 3207 6702
rect 10501 6762 10567 6765
rect 33317 6762 33383 6765
rect 10501 6760 33383 6762
rect 10501 6704 10506 6760
rect 10562 6704 33322 6760
rect 33378 6704 33383 6760
rect 10501 6702 33383 6704
rect 10501 6699 10567 6702
rect 33317 6699 33383 6702
rect 2865 6626 2931 6629
rect 7005 6626 7071 6629
rect 2865 6624 7071 6626
rect 2865 6568 2870 6624
rect 2926 6568 7010 6624
rect 7066 6568 7071 6624
rect 2865 6566 7071 6568
rect 2865 6563 2931 6566
rect 7005 6563 7071 6566
rect 10869 6626 10935 6629
rect 13486 6626 13492 6628
rect 10869 6624 13492 6626
rect 10869 6568 10874 6624
rect 10930 6568 13492 6624
rect 10869 6566 13492 6568
rect 10869 6563 10935 6566
rect 13486 6564 13492 6566
rect 13556 6564 13562 6628
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 4245 6490 4311 6493
rect 0 6488 4311 6490
rect 0 6432 4250 6488
rect 4306 6432 4311 6488
rect 0 6430 4311 6432
rect 0 6400 800 6430
rect 4245 6427 4311 6430
rect 6913 6490 6979 6493
rect 7598 6490 7604 6492
rect 6913 6488 7604 6490
rect 6913 6432 6918 6488
rect 6974 6432 7604 6488
rect 6913 6430 7604 6432
rect 6913 6427 6979 6430
rect 7598 6428 7604 6430
rect 7668 6428 7674 6492
rect 8477 6490 8543 6493
rect 17166 6490 17172 6492
rect 8477 6488 17172 6490
rect 8477 6432 8482 6488
rect 8538 6432 17172 6488
rect 8477 6430 17172 6432
rect 8477 6427 8543 6430
rect 17166 6428 17172 6430
rect 17236 6428 17242 6492
rect 3141 6354 3207 6357
rect 3969 6354 4035 6357
rect 3141 6352 4035 6354
rect 3141 6296 3146 6352
rect 3202 6296 3974 6352
rect 4030 6296 4035 6352
rect 3141 6294 4035 6296
rect 3141 6291 3207 6294
rect 3969 6291 4035 6294
rect 4153 6354 4219 6357
rect 24710 6354 24716 6356
rect 4153 6352 24716 6354
rect 4153 6296 4158 6352
rect 4214 6296 24716 6352
rect 4153 6294 24716 6296
rect 4153 6291 4219 6294
rect 24710 6292 24716 6294
rect 24780 6292 24786 6356
rect 2865 6218 2931 6221
rect 13537 6218 13603 6221
rect 2865 6216 13603 6218
rect 2865 6160 2870 6216
rect 2926 6160 13542 6216
rect 13598 6160 13603 6216
rect 2865 6158 13603 6160
rect 2865 6155 2931 6158
rect 13537 6155 13603 6158
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 4153 6082 4219 6085
rect 4286 6082 4292 6084
rect 4153 6080 4292 6082
rect 4153 6024 4158 6080
rect 4214 6024 4292 6080
rect 4153 6022 4292 6024
rect 4153 6019 4219 6022
rect 4286 6020 4292 6022
rect 4356 6020 4362 6084
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 4153 5810 4219 5813
rect 22686 5810 22692 5812
rect 4153 5808 22692 5810
rect 4153 5752 4158 5808
rect 4214 5752 22692 5808
rect 4153 5750 22692 5752
rect 4153 5747 4219 5750
rect 22686 5748 22692 5750
rect 22756 5748 22762 5812
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 7833 5674 7899 5677
rect 16614 5674 16620 5676
rect 7833 5672 16620 5674
rect 7833 5616 7838 5672
rect 7894 5616 16620 5672
rect 7833 5614 16620 5616
rect 7833 5611 7899 5614
rect 16614 5612 16620 5614
rect 16684 5612 16690 5676
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1577 4858 1643 4861
rect 0 4856 1643 4858
rect 0 4800 1582 4856
rect 1638 4800 1643 4856
rect 0 4798 1643 4800
rect 0 4768 800 4798
rect 1577 4795 1643 4798
rect 3325 4722 3391 4725
rect 8293 4722 8359 4725
rect 3325 4720 8359 4722
rect 3325 4664 3330 4720
rect 3386 4664 8298 4720
rect 8354 4664 8359 4720
rect 3325 4662 8359 4664
rect 3325 4659 3391 4662
rect 8293 4659 8359 4662
rect 0 4450 800 4480
rect 3693 4450 3759 4453
rect 0 4448 3759 4450
rect 0 4392 3698 4448
rect 3754 4392 3759 4448
rect 0 4390 3759 4392
rect 0 4360 800 4390
rect 3693 4387 3759 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 1209 4042 1275 4045
rect 0 4040 1275 4042
rect 0 3984 1214 4040
rect 1270 3984 1275 4040
rect 0 3982 1275 3984
rect 0 3952 800 3982
rect 1209 3979 1275 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 4061 3226 4127 3229
rect 0 3224 4127 3226
rect 0 3168 4066 3224
rect 4122 3168 4127 3224
rect 0 3166 4127 3168
rect 0 3136 800 3166
rect 4061 3163 4127 3166
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
<< via3 >>
rect 12572 26284 12636 26348
rect 33364 26012 33428 26076
rect 12756 25876 12820 25940
rect 11468 25740 11532 25804
rect 16620 25468 16684 25532
rect 14412 25332 14476 25396
rect 24900 25196 24964 25260
rect 14228 25060 14292 25124
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 15700 24380 15764 24444
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 13676 23700 13740 23764
rect 15148 23564 15212 23628
rect 19932 23564 19996 23628
rect 9628 23428 9692 23492
rect 15332 23488 15396 23492
rect 15332 23432 15346 23488
rect 15346 23432 15396 23488
rect 15332 23428 15396 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 11468 22884 11532 22948
rect 13860 23020 13924 23084
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 11652 22748 11716 22812
rect 12572 22748 12636 22812
rect 3556 22612 3620 22676
rect 24716 22672 24780 22676
rect 24716 22616 24730 22672
rect 24730 22616 24780 22672
rect 24716 22612 24780 22616
rect 4660 22400 4724 22404
rect 4660 22344 4674 22400
rect 4674 22344 4724 22400
rect 4660 22340 4724 22344
rect 7420 22400 7484 22404
rect 7420 22344 7434 22400
rect 7434 22344 7484 22400
rect 7420 22340 7484 22344
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 19564 22264 19628 22268
rect 19564 22208 19614 22264
rect 19614 22208 19628 22264
rect 19564 22204 19628 22208
rect 2636 21796 2700 21860
rect 14228 21932 14292 21996
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2452 21660 2516 21724
rect 33364 21720 33428 21724
rect 33364 21664 33414 21720
rect 33414 21664 33428 21720
rect 33364 21660 33428 21664
rect 10732 21388 10796 21452
rect 11100 21312 11164 21316
rect 11100 21256 11150 21312
rect 11150 21256 11164 21312
rect 11100 21252 11164 21256
rect 13676 21252 13740 21316
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 19748 21116 19812 21180
rect 6684 20980 6748 21044
rect 10916 20980 10980 21044
rect 14044 20708 14108 20772
rect 14412 20708 14476 20772
rect 22692 20708 22756 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 5764 20572 5828 20636
rect 10364 20572 10428 20636
rect 18644 20572 18708 20636
rect 19380 20436 19444 20500
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 1164 19756 1228 19820
rect 5580 19484 5644 19548
rect 3740 19348 3804 19412
rect 6132 19348 6196 19412
rect 12756 19620 12820 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 22508 19544 22572 19548
rect 22508 19488 22522 19544
rect 22522 19488 22572 19544
rect 22508 19484 22572 19488
rect 8708 19348 8772 19412
rect 10180 19272 10244 19276
rect 10180 19216 10194 19272
rect 10194 19216 10244 19272
rect 10180 19212 10244 19216
rect 11284 19348 11348 19412
rect 17172 19348 17236 19412
rect 15516 19076 15580 19140
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 24900 18940 24964 19004
rect 8340 18728 8404 18732
rect 8340 18672 8354 18728
rect 8354 18672 8404 18728
rect 8340 18668 8404 18672
rect 1348 18532 1412 18596
rect 7236 18592 7300 18596
rect 7236 18536 7286 18592
rect 7286 18536 7300 18592
rect 7236 18532 7300 18536
rect 9812 18592 9876 18596
rect 9812 18536 9826 18592
rect 9826 18536 9876 18592
rect 9812 18532 9876 18536
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 980 18396 1044 18460
rect 12020 18532 12084 18596
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 11836 18456 11900 18460
rect 11836 18400 11850 18456
rect 11850 18400 11900 18456
rect 11836 18396 11900 18400
rect 12204 18396 12268 18460
rect 9996 18260 10060 18324
rect 15516 18260 15580 18324
rect 8524 18184 8588 18188
rect 8524 18128 8574 18184
rect 8574 18128 8588 18184
rect 8524 18124 8588 18128
rect 4108 17988 4172 18052
rect 16252 18048 16316 18052
rect 16252 17992 16302 18048
rect 16302 17992 16316 18048
rect 16252 17988 16316 17992
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 4476 17852 4540 17916
rect 18460 18048 18524 18052
rect 18460 17992 18474 18048
rect 18474 17992 18524 18048
rect 18460 17988 18524 17992
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 3924 17580 3988 17644
rect 16252 17580 16316 17644
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 9444 17308 9508 17372
rect 9812 17308 9876 17372
rect 1532 17172 1596 17236
rect 3556 17172 3620 17236
rect 5028 17036 5092 17100
rect 14780 17036 14844 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 9260 16764 9324 16828
rect 12204 16764 12268 16828
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 13860 16356 13924 16420
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 12020 16220 12084 16284
rect 8524 15872 8588 15876
rect 8524 15816 8538 15872
rect 8538 15816 8588 15872
rect 8524 15812 8588 15816
rect 8892 15812 8956 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 19380 15812 19444 15876
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 11284 15404 11348 15468
rect 4292 15328 4356 15332
rect 4292 15272 4342 15328
rect 4342 15272 4356 15328
rect 4292 15268 4356 15272
rect 13492 15328 13556 15332
rect 13492 15272 13542 15328
rect 13542 15272 13556 15328
rect 13492 15268 13556 15272
rect 14964 15328 15028 15332
rect 14964 15272 15014 15328
rect 15014 15272 15028 15328
rect 14964 15268 15028 15272
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 9076 15132 9140 15196
rect 3740 14860 3804 14924
rect 5580 14724 5644 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 8892 14588 8956 14652
rect 7604 14316 7668 14380
rect 8892 14376 8956 14380
rect 8892 14320 8906 14376
rect 8906 14320 8956 14376
rect 8892 14316 8956 14320
rect 8340 14180 8404 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 5580 13832 5644 13836
rect 5580 13776 5594 13832
rect 5594 13776 5644 13832
rect 5580 13772 5644 13776
rect 5028 13636 5092 13700
rect 5212 13696 5276 13700
rect 5212 13640 5262 13696
rect 5262 13640 5276 13696
rect 5212 13636 5276 13640
rect 12204 13636 12268 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 3372 13500 3436 13564
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 1900 13364 1964 13428
rect 14780 13364 14844 13428
rect 18644 13364 18708 13428
rect 19748 13364 19812 13428
rect 10916 13228 10980 13292
rect 9996 13092 10060 13156
rect 19932 13092 19996 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 9260 12956 9324 13020
rect 12756 13016 12820 13020
rect 12756 12960 12770 13016
rect 12770 12960 12820 13016
rect 12756 12956 12820 12960
rect 13676 12956 13740 13020
rect 5948 12820 6012 12884
rect 19564 12820 19628 12884
rect 9996 12684 10060 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 4292 12336 4356 12340
rect 4292 12280 4342 12336
rect 4342 12280 4356 12336
rect 4292 12276 4356 12280
rect 8708 12140 8772 12204
rect 4292 12004 4356 12068
rect 16252 12064 16316 12068
rect 16252 12008 16302 12064
rect 16302 12008 16316 12064
rect 16252 12004 16316 12008
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2452 11928 2516 11932
rect 2452 11872 2466 11928
rect 2466 11872 2516 11928
rect 2452 11868 2516 11872
rect 3740 11732 3804 11796
rect 5396 11732 5460 11796
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 4660 11324 4724 11388
rect 13676 11324 13740 11388
rect 14228 11384 14292 11388
rect 14228 11328 14242 11384
rect 14242 11328 14292 11384
rect 14228 11324 14292 11328
rect 9996 11052 10060 11116
rect 18460 11188 18524 11252
rect 1900 10976 1964 10980
rect 1900 10920 1914 10976
rect 1914 10920 1964 10976
rect 1900 10916 1964 10920
rect 7236 10916 7300 10980
rect 9812 10976 9876 10980
rect 9812 10920 9826 10976
rect 9826 10920 9876 10976
rect 9812 10916 9876 10920
rect 12572 10916 12636 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 3924 10780 3988 10844
rect 1348 10644 1412 10708
rect 5948 10644 6012 10708
rect 11836 10644 11900 10708
rect 2636 10372 2700 10436
rect 9260 10372 9324 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 15332 10100 15396 10164
rect 3556 9964 3620 10028
rect 4476 9888 4540 9892
rect 4476 9832 4526 9888
rect 4526 9832 4540 9888
rect 4476 9828 4540 9832
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 5764 9752 5828 9756
rect 5764 9696 5814 9752
rect 5814 9696 5828 9752
rect 5764 9692 5828 9696
rect 6132 9692 6196 9756
rect 6684 9692 6748 9756
rect 1532 9616 1596 9620
rect 1532 9560 1546 9616
rect 1546 9560 1596 9616
rect 1532 9556 1596 9560
rect 3372 9616 3436 9620
rect 3372 9560 3386 9616
rect 3386 9560 3436 9616
rect 3372 9556 3436 9560
rect 4108 9556 4172 9620
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 10732 9752 10796 9756
rect 10732 9696 10746 9752
rect 10746 9696 10796 9752
rect 10732 9692 10796 9696
rect 12756 9692 12820 9756
rect 14964 9692 15028 9756
rect 14044 9556 14108 9620
rect 15148 9556 15212 9620
rect 980 9420 1044 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 12756 9148 12820 9212
rect 3740 9012 3804 9076
rect 5396 9012 5460 9076
rect 9444 9012 9508 9076
rect 10364 9012 10428 9076
rect 15148 8740 15212 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 11100 8664 11164 8668
rect 11100 8608 11114 8664
rect 11114 8608 11164 8664
rect 11100 8604 11164 8608
rect 11468 8604 11532 8668
rect 11652 8664 11716 8668
rect 11652 8608 11666 8664
rect 11666 8608 11716 8664
rect 11652 8604 11716 8608
rect 9076 8468 9140 8532
rect 15516 8468 15580 8532
rect 5212 8196 5276 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 12204 8060 12268 8124
rect 15700 7652 15764 7716
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 1164 7516 1228 7580
rect 3556 7380 3620 7444
rect 7420 7440 7484 7444
rect 7420 7384 7434 7440
rect 7434 7384 7484 7440
rect 7420 7380 7484 7384
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 13676 7108 13740 7172
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 10180 6972 10244 7036
rect 8892 6836 8956 6900
rect 22508 6972 22572 7036
rect 13492 6564 13556 6628
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 7604 6428 7668 6492
rect 17172 6428 17236 6492
rect 24716 6292 24780 6356
rect 4292 6020 4356 6084
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 22692 5748 22756 5812
rect 16620 5612 16684 5676
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 12571 26348 12637 26349
rect 12571 26284 12572 26348
rect 12636 26284 12637 26348
rect 12571 26283 12637 26284
rect 11467 25804 11533 25805
rect 11467 25740 11468 25804
rect 11532 25740 11533 25804
rect 11467 25739 11533 25740
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 9627 23492 9693 23493
rect 9627 23428 9628 23492
rect 9692 23428 9693 23492
rect 9627 23427 9693 23428
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 3555 22676 3621 22677
rect 3555 22612 3556 22676
rect 3620 22612 3621 22676
rect 3555 22611 3621 22612
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2635 21860 2701 21861
rect 2635 21796 2636 21860
rect 2700 21796 2701 21860
rect 2635 21795 2701 21796
rect 2451 21724 2517 21725
rect 2451 21660 2452 21724
rect 2516 21660 2517 21724
rect 2451 21659 2517 21660
rect 1163 19820 1229 19821
rect 1163 19756 1164 19820
rect 1228 19756 1229 19820
rect 1163 19755 1229 19756
rect 979 18460 1045 18461
rect 979 18396 980 18460
rect 1044 18396 1045 18460
rect 979 18395 1045 18396
rect 982 9485 1042 18395
rect 979 9484 1045 9485
rect 979 9420 980 9484
rect 1044 9420 1045 9484
rect 979 9419 1045 9420
rect 1166 7581 1226 19755
rect 1347 18596 1413 18597
rect 1347 18532 1348 18596
rect 1412 18532 1413 18596
rect 1347 18531 1413 18532
rect 1350 10709 1410 18531
rect 1531 17236 1597 17237
rect 1531 17172 1532 17236
rect 1596 17172 1597 17236
rect 1531 17171 1597 17172
rect 1347 10708 1413 10709
rect 1347 10644 1348 10708
rect 1412 10644 1413 10708
rect 1347 10643 1413 10644
rect 1534 9621 1594 17171
rect 1899 13428 1965 13429
rect 1899 13364 1900 13428
rect 1964 13364 1965 13428
rect 1899 13363 1965 13364
rect 1902 10981 1962 13363
rect 2454 11933 2514 21659
rect 2451 11932 2517 11933
rect 2451 11868 2452 11932
rect 2516 11868 2517 11932
rect 2451 11867 2517 11868
rect 1899 10980 1965 10981
rect 1899 10916 1900 10980
rect 1964 10916 1965 10980
rect 1899 10915 1965 10916
rect 2638 10437 2698 21795
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 3558 17237 3618 22611
rect 4659 22404 4725 22405
rect 4659 22340 4660 22404
rect 4724 22340 4725 22404
rect 4659 22339 4725 22340
rect 7419 22404 7485 22405
rect 7419 22340 7420 22404
rect 7484 22340 7485 22404
rect 7419 22339 7485 22340
rect 3739 19412 3805 19413
rect 3739 19348 3740 19412
rect 3804 19348 3805 19412
rect 3739 19347 3805 19348
rect 3555 17236 3621 17237
rect 3555 17172 3556 17236
rect 3620 17172 3621 17236
rect 3555 17171 3621 17172
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 3742 14925 3802 19347
rect 4107 18052 4173 18053
rect 4107 17988 4108 18052
rect 4172 17988 4173 18052
rect 4107 17987 4173 17988
rect 3923 17644 3989 17645
rect 3923 17580 3924 17644
rect 3988 17580 3989 17644
rect 3923 17579 3989 17580
rect 3739 14924 3805 14925
rect 3739 14860 3740 14924
rect 3804 14860 3805 14924
rect 3739 14859 3805 14860
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 3371 13564 3437 13565
rect 3371 13500 3372 13564
rect 3436 13500 3437 13564
rect 3371 13499 3437 13500
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2635 10436 2701 10437
rect 2635 10372 2636 10436
rect 2700 10372 2701 10436
rect 2635 10371 2701 10372
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 1531 9620 1597 9621
rect 1531 9556 1532 9620
rect 1596 9556 1597 9620
rect 1531 9555 1597 9556
rect 2944 9280 3264 10304
rect 3374 9621 3434 13499
rect 3739 11796 3805 11797
rect 3739 11732 3740 11796
rect 3804 11732 3805 11796
rect 3739 11731 3805 11732
rect 3555 10028 3621 10029
rect 3555 9964 3556 10028
rect 3620 9964 3621 10028
rect 3555 9963 3621 9964
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 1163 7580 1229 7581
rect 1163 7516 1164 7580
rect 1228 7516 1229 7580
rect 1163 7515 1229 7516
rect 2944 7104 3264 8128
rect 3558 7445 3618 9963
rect 3742 9077 3802 11731
rect 3926 10845 3986 17579
rect 3923 10844 3989 10845
rect 3923 10780 3924 10844
rect 3988 10780 3989 10844
rect 3923 10779 3989 10780
rect 4110 9621 4170 17987
rect 4475 17916 4541 17917
rect 4475 17852 4476 17916
rect 4540 17852 4541 17916
rect 4475 17851 4541 17852
rect 4291 15332 4357 15333
rect 4291 15268 4292 15332
rect 4356 15268 4357 15332
rect 4291 15267 4357 15268
rect 4294 12341 4354 15267
rect 4291 12340 4357 12341
rect 4291 12276 4292 12340
rect 4356 12276 4357 12340
rect 4291 12275 4357 12276
rect 4291 12068 4357 12069
rect 4291 12004 4292 12068
rect 4356 12004 4357 12068
rect 4291 12003 4357 12004
rect 4107 9620 4173 9621
rect 4107 9556 4108 9620
rect 4172 9556 4173 9620
rect 4107 9555 4173 9556
rect 3739 9076 3805 9077
rect 3739 9012 3740 9076
rect 3804 9012 3805 9076
rect 3739 9011 3805 9012
rect 3555 7444 3621 7445
rect 3555 7380 3556 7444
rect 3620 7380 3621 7444
rect 3555 7379 3621 7380
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 4294 6085 4354 12003
rect 4478 9893 4538 17851
rect 4662 11389 4722 22339
rect 6683 21044 6749 21045
rect 6683 20980 6684 21044
rect 6748 20980 6749 21044
rect 6683 20979 6749 20980
rect 5763 20636 5829 20637
rect 5763 20572 5764 20636
rect 5828 20572 5829 20636
rect 5763 20571 5829 20572
rect 5579 19548 5645 19549
rect 5579 19484 5580 19548
rect 5644 19484 5645 19548
rect 5579 19483 5645 19484
rect 5027 17100 5093 17101
rect 5027 17036 5028 17100
rect 5092 17036 5093 17100
rect 5027 17035 5093 17036
rect 5030 13701 5090 17035
rect 5582 14789 5642 19483
rect 5579 14788 5645 14789
rect 5579 14724 5580 14788
rect 5644 14724 5645 14788
rect 5579 14723 5645 14724
rect 5582 13837 5642 14723
rect 5579 13836 5645 13837
rect 5579 13772 5580 13836
rect 5644 13772 5645 13836
rect 5579 13771 5645 13772
rect 5027 13700 5093 13701
rect 5027 13636 5028 13700
rect 5092 13636 5093 13700
rect 5027 13635 5093 13636
rect 5211 13700 5277 13701
rect 5211 13636 5212 13700
rect 5276 13636 5277 13700
rect 5211 13635 5277 13636
rect 4659 11388 4725 11389
rect 4659 11324 4660 11388
rect 4724 11324 4725 11388
rect 4659 11323 4725 11324
rect 4475 9892 4541 9893
rect 4475 9828 4476 9892
rect 4540 9828 4541 9892
rect 4475 9827 4541 9828
rect 5214 8261 5274 13635
rect 5395 11796 5461 11797
rect 5395 11732 5396 11796
rect 5460 11732 5461 11796
rect 5395 11731 5461 11732
rect 5398 9077 5458 11731
rect 5766 9757 5826 20571
rect 6131 19412 6197 19413
rect 6131 19348 6132 19412
rect 6196 19348 6197 19412
rect 6131 19347 6197 19348
rect 5947 12884 6013 12885
rect 5947 12820 5948 12884
rect 6012 12820 6013 12884
rect 5947 12819 6013 12820
rect 5950 10709 6010 12819
rect 5947 10708 6013 10709
rect 5947 10644 5948 10708
rect 6012 10644 6013 10708
rect 5947 10643 6013 10644
rect 6134 9757 6194 19347
rect 6686 9757 6746 20979
rect 7235 18596 7301 18597
rect 7235 18532 7236 18596
rect 7300 18532 7301 18596
rect 7235 18531 7301 18532
rect 7238 10981 7298 18531
rect 7235 10980 7301 10981
rect 7235 10916 7236 10980
rect 7300 10916 7301 10980
rect 7235 10915 7301 10916
rect 5763 9756 5829 9757
rect 5763 9692 5764 9756
rect 5828 9692 5829 9756
rect 5763 9691 5829 9692
rect 6131 9756 6197 9757
rect 6131 9692 6132 9756
rect 6196 9692 6197 9756
rect 6131 9691 6197 9692
rect 6683 9756 6749 9757
rect 6683 9692 6684 9756
rect 6748 9692 6749 9756
rect 6683 9691 6749 9692
rect 5395 9076 5461 9077
rect 5395 9012 5396 9076
rect 5460 9012 5461 9076
rect 5395 9011 5461 9012
rect 5211 8260 5277 8261
rect 5211 8196 5212 8260
rect 5276 8196 5277 8260
rect 5211 8195 5277 8196
rect 7422 7445 7482 22339
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 8707 19412 8773 19413
rect 8707 19348 8708 19412
rect 8772 19348 8773 19412
rect 8707 19347 8773 19348
rect 8339 18732 8405 18733
rect 8339 18668 8340 18732
rect 8404 18668 8405 18732
rect 8339 18667 8405 18668
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7603 14380 7669 14381
rect 7603 14316 7604 14380
rect 7668 14316 7669 14380
rect 7603 14315 7669 14316
rect 7419 7444 7485 7445
rect 7419 7380 7420 7444
rect 7484 7380 7485 7444
rect 7419 7379 7485 7380
rect 7606 6493 7666 14315
rect 7944 14176 8264 15200
rect 8342 14245 8402 18667
rect 8523 18188 8589 18189
rect 8523 18124 8524 18188
rect 8588 18124 8589 18188
rect 8523 18123 8589 18124
rect 8526 15877 8586 18123
rect 8523 15876 8589 15877
rect 8523 15812 8524 15876
rect 8588 15812 8589 15876
rect 8523 15811 8589 15812
rect 8339 14244 8405 14245
rect 8339 14180 8340 14244
rect 8404 14180 8405 14244
rect 8339 14179 8405 14180
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 8710 12205 8770 19347
rect 9443 17372 9509 17373
rect 9443 17308 9444 17372
rect 9508 17308 9509 17372
rect 9443 17307 9509 17308
rect 9259 16828 9325 16829
rect 9259 16764 9260 16828
rect 9324 16764 9325 16828
rect 9259 16763 9325 16764
rect 8891 15876 8957 15877
rect 8891 15812 8892 15876
rect 8956 15812 8957 15876
rect 8891 15811 8957 15812
rect 8894 14653 8954 15811
rect 9075 15196 9141 15197
rect 9075 15132 9076 15196
rect 9140 15132 9141 15196
rect 9075 15131 9141 15132
rect 8891 14652 8957 14653
rect 8891 14588 8892 14652
rect 8956 14588 8957 14652
rect 8891 14587 8957 14588
rect 8891 14380 8957 14381
rect 8891 14316 8892 14380
rect 8956 14316 8957 14380
rect 8891 14315 8957 14316
rect 8707 12204 8773 12205
rect 8707 12140 8708 12204
rect 8772 12140 8773 12204
rect 8707 12139 8773 12140
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 8894 6901 8954 14315
rect 9078 8533 9138 15131
rect 9262 13021 9322 16763
rect 9259 13020 9325 13021
rect 9259 12956 9260 13020
rect 9324 12956 9325 13020
rect 9259 12955 9325 12956
rect 9262 10437 9322 12955
rect 9259 10436 9325 10437
rect 9259 10372 9260 10436
rect 9324 10372 9325 10436
rect 9259 10371 9325 10372
rect 9446 9077 9506 17307
rect 9630 14650 9690 23427
rect 11470 22949 11530 25739
rect 11467 22948 11533 22949
rect 11467 22884 11468 22948
rect 11532 22884 11533 22948
rect 11467 22883 11533 22884
rect 10731 21452 10797 21453
rect 10731 21388 10732 21452
rect 10796 21388 10797 21452
rect 10731 21387 10797 21388
rect 10363 20636 10429 20637
rect 10363 20572 10364 20636
rect 10428 20572 10429 20636
rect 10363 20571 10429 20572
rect 10179 19276 10245 19277
rect 10179 19212 10180 19276
rect 10244 19212 10245 19276
rect 10179 19211 10245 19212
rect 9811 18596 9877 18597
rect 9811 18532 9812 18596
rect 9876 18532 9877 18596
rect 9811 18531 9877 18532
rect 9814 17373 9874 18531
rect 9995 18324 10061 18325
rect 9995 18260 9996 18324
rect 10060 18260 10061 18324
rect 9995 18259 10061 18260
rect 9811 17372 9877 17373
rect 9811 17308 9812 17372
rect 9876 17308 9877 17372
rect 9811 17307 9877 17308
rect 9630 14590 9874 14650
rect 9814 10981 9874 14590
rect 9998 13157 10058 18259
rect 9995 13156 10061 13157
rect 9995 13092 9996 13156
rect 10060 13092 10061 13156
rect 9995 13091 10061 13092
rect 9995 12748 10061 12749
rect 9995 12684 9996 12748
rect 10060 12684 10061 12748
rect 9995 12683 10061 12684
rect 9998 11117 10058 12683
rect 9995 11116 10061 11117
rect 9995 11052 9996 11116
rect 10060 11052 10061 11116
rect 9995 11051 10061 11052
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 9443 9076 9509 9077
rect 9443 9012 9444 9076
rect 9508 9012 9509 9076
rect 9443 9011 9509 9012
rect 9075 8532 9141 8533
rect 9075 8468 9076 8532
rect 9140 8468 9141 8532
rect 9075 8467 9141 8468
rect 10182 7037 10242 19211
rect 10366 9077 10426 20571
rect 10734 9757 10794 21387
rect 11099 21316 11165 21317
rect 11099 21252 11100 21316
rect 11164 21252 11165 21316
rect 11099 21251 11165 21252
rect 10915 21044 10981 21045
rect 10915 20980 10916 21044
rect 10980 20980 10981 21044
rect 10915 20979 10981 20980
rect 10918 13293 10978 20979
rect 10915 13292 10981 13293
rect 10915 13228 10916 13292
rect 10980 13228 10981 13292
rect 10915 13227 10981 13228
rect 10731 9756 10797 9757
rect 10731 9692 10732 9756
rect 10796 9692 10797 9756
rect 10731 9691 10797 9692
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 11102 8669 11162 21251
rect 11283 19412 11349 19413
rect 11283 19348 11284 19412
rect 11348 19348 11349 19412
rect 11283 19347 11349 19348
rect 11286 15469 11346 19347
rect 11283 15468 11349 15469
rect 11283 15404 11284 15468
rect 11348 15404 11349 15468
rect 11283 15403 11349 15404
rect 11470 8669 11530 22883
rect 12574 22813 12634 26283
rect 33363 26076 33429 26077
rect 33363 26012 33364 26076
rect 33428 26012 33429 26076
rect 33363 26011 33429 26012
rect 12755 25940 12821 25941
rect 12755 25876 12756 25940
rect 12820 25876 12821 25940
rect 12755 25875 12821 25876
rect 11651 22812 11717 22813
rect 11651 22748 11652 22812
rect 11716 22748 11717 22812
rect 11651 22747 11717 22748
rect 12571 22812 12637 22813
rect 12571 22748 12572 22812
rect 12636 22748 12637 22812
rect 12571 22747 12637 22748
rect 11654 8669 11714 22747
rect 12574 22110 12634 22747
rect 12390 22050 12634 22110
rect 12390 21450 12450 22050
rect 12390 21390 12634 21450
rect 12019 18596 12085 18597
rect 12019 18532 12020 18596
rect 12084 18532 12085 18596
rect 12019 18531 12085 18532
rect 11835 18460 11901 18461
rect 11835 18396 11836 18460
rect 11900 18396 11901 18460
rect 11835 18395 11901 18396
rect 11838 10709 11898 18395
rect 12022 16285 12082 18531
rect 12203 18460 12269 18461
rect 12203 18396 12204 18460
rect 12268 18396 12269 18460
rect 12203 18395 12269 18396
rect 12206 16829 12266 18395
rect 12203 16828 12269 16829
rect 12203 16764 12204 16828
rect 12268 16764 12269 16828
rect 12203 16763 12269 16764
rect 12019 16284 12085 16285
rect 12019 16220 12020 16284
rect 12084 16220 12085 16284
rect 12019 16219 12085 16220
rect 12203 13700 12269 13701
rect 12203 13636 12204 13700
rect 12268 13636 12269 13700
rect 12203 13635 12269 13636
rect 11835 10708 11901 10709
rect 11835 10644 11836 10708
rect 11900 10644 11901 10708
rect 11835 10643 11901 10644
rect 11099 8668 11165 8669
rect 11099 8604 11100 8668
rect 11164 8604 11165 8668
rect 11099 8603 11165 8604
rect 11467 8668 11533 8669
rect 11467 8604 11468 8668
rect 11532 8604 11533 8668
rect 11467 8603 11533 8604
rect 11651 8668 11717 8669
rect 11651 8604 11652 8668
rect 11716 8604 11717 8668
rect 11651 8603 11717 8604
rect 12206 8125 12266 13635
rect 12574 10981 12634 21390
rect 12758 19685 12818 25875
rect 16619 25532 16685 25533
rect 16619 25468 16620 25532
rect 16684 25468 16685 25532
rect 16619 25467 16685 25468
rect 14411 25396 14477 25397
rect 14411 25332 14412 25396
rect 14476 25332 14477 25396
rect 14411 25331 14477 25332
rect 14227 25124 14293 25125
rect 14227 25060 14228 25124
rect 14292 25060 14293 25124
rect 14227 25059 14293 25060
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 13675 23764 13741 23765
rect 13675 23700 13676 23764
rect 13740 23700 13741 23764
rect 13675 23699 13741 23700
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 13678 21317 13738 23699
rect 13859 23084 13925 23085
rect 13859 23020 13860 23084
rect 13924 23020 13925 23084
rect 13859 23019 13925 23020
rect 13675 21316 13741 21317
rect 13675 21252 13676 21316
rect 13740 21252 13741 21316
rect 13675 21251 13741 21252
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12755 19684 12821 19685
rect 12755 19620 12756 19684
rect 12820 19620 12821 19684
rect 12755 19619 12821 19620
rect 12758 13021 12818 19619
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 13491 15332 13557 15333
rect 13491 15268 13492 15332
rect 13556 15268 13557 15332
rect 13491 15267 13557 15268
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12755 13020 12821 13021
rect 12755 12956 12756 13020
rect 12820 12956 12821 13020
rect 12755 12955 12821 12956
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12571 10980 12637 10981
rect 12571 10916 12572 10980
rect 12636 10916 12637 10980
rect 12571 10915 12637 10916
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12755 9756 12821 9757
rect 12755 9692 12756 9756
rect 12820 9692 12821 9756
rect 12755 9691 12821 9692
rect 12758 9213 12818 9691
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12755 9212 12821 9213
rect 12755 9148 12756 9212
rect 12820 9148 12821 9212
rect 12755 9147 12821 9148
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12203 8124 12269 8125
rect 12203 8060 12204 8124
rect 12268 8060 12269 8124
rect 12203 8059 12269 8060
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 10179 7036 10245 7037
rect 10179 6972 10180 7036
rect 10244 6972 10245 7036
rect 10179 6971 10245 6972
rect 8891 6900 8957 6901
rect 8891 6836 8892 6900
rect 8956 6836 8957 6900
rect 8891 6835 8957 6836
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7603 6492 7669 6493
rect 7603 6428 7604 6492
rect 7668 6428 7669 6492
rect 7603 6427 7669 6428
rect 4291 6084 4357 6085
rect 4291 6020 4292 6084
rect 4356 6020 4357 6084
rect 4291 6019 4357 6020
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 6016 13264 7040
rect 13494 6629 13554 15267
rect 13678 13021 13738 21251
rect 13862 16421 13922 23019
rect 14230 21997 14290 25059
rect 14227 21996 14293 21997
rect 14227 21932 14228 21996
rect 14292 21932 14293 21996
rect 14227 21931 14293 21932
rect 14043 20772 14109 20773
rect 14043 20708 14044 20772
rect 14108 20708 14109 20772
rect 14043 20707 14109 20708
rect 13859 16420 13925 16421
rect 13859 16356 13860 16420
rect 13924 16356 13925 16420
rect 13859 16355 13925 16356
rect 13675 13020 13741 13021
rect 13675 12956 13676 13020
rect 13740 12956 13741 13020
rect 13675 12955 13741 12956
rect 13675 11388 13741 11389
rect 13675 11324 13676 11388
rect 13740 11324 13741 11388
rect 13675 11323 13741 11324
rect 13678 7173 13738 11323
rect 14046 9621 14106 20707
rect 14230 11389 14290 21931
rect 14414 20773 14474 25331
rect 15699 24444 15765 24445
rect 15699 24380 15700 24444
rect 15764 24380 15765 24444
rect 15699 24379 15765 24380
rect 15147 23628 15213 23629
rect 15147 23564 15148 23628
rect 15212 23564 15213 23628
rect 15147 23563 15213 23564
rect 14411 20772 14477 20773
rect 14411 20708 14412 20772
rect 14476 20708 14477 20772
rect 14411 20707 14477 20708
rect 14779 17100 14845 17101
rect 14779 17036 14780 17100
rect 14844 17036 14845 17100
rect 14779 17035 14845 17036
rect 14782 13429 14842 17035
rect 14963 15332 15029 15333
rect 14963 15268 14964 15332
rect 15028 15268 15029 15332
rect 14963 15267 15029 15268
rect 14779 13428 14845 13429
rect 14779 13364 14780 13428
rect 14844 13364 14845 13428
rect 14779 13363 14845 13364
rect 14227 11388 14293 11389
rect 14227 11324 14228 11388
rect 14292 11324 14293 11388
rect 14227 11323 14293 11324
rect 14966 9757 15026 15267
rect 14963 9756 15029 9757
rect 14963 9692 14964 9756
rect 15028 9692 15029 9756
rect 14963 9691 15029 9692
rect 15150 9621 15210 23563
rect 15331 23492 15397 23493
rect 15331 23428 15332 23492
rect 15396 23428 15397 23492
rect 15331 23427 15397 23428
rect 15334 10165 15394 23427
rect 15515 19140 15581 19141
rect 15515 19076 15516 19140
rect 15580 19076 15581 19140
rect 15515 19075 15581 19076
rect 15518 18325 15578 19075
rect 15515 18324 15581 18325
rect 15515 18260 15516 18324
rect 15580 18260 15581 18324
rect 15515 18259 15581 18260
rect 15331 10164 15397 10165
rect 15331 10100 15332 10164
rect 15396 10100 15397 10164
rect 15331 10099 15397 10100
rect 14043 9620 14109 9621
rect 14043 9556 14044 9620
rect 14108 9556 14109 9620
rect 14043 9555 14109 9556
rect 15147 9620 15213 9621
rect 15147 9556 15148 9620
rect 15212 9556 15213 9620
rect 15147 9555 15213 9556
rect 15150 8805 15210 9555
rect 15147 8804 15213 8805
rect 15147 8740 15148 8804
rect 15212 8740 15213 8804
rect 15147 8739 15213 8740
rect 15518 8533 15578 18259
rect 15515 8532 15581 8533
rect 15515 8468 15516 8532
rect 15580 8468 15581 8532
rect 15515 8467 15581 8468
rect 15702 7717 15762 24379
rect 16251 18052 16317 18053
rect 16251 17988 16252 18052
rect 16316 17988 16317 18052
rect 16251 17987 16317 17988
rect 16254 17645 16314 17987
rect 16251 17644 16317 17645
rect 16251 17580 16252 17644
rect 16316 17580 16317 17644
rect 16251 17579 16317 17580
rect 16254 12069 16314 17579
rect 16251 12068 16317 12069
rect 16251 12004 16252 12068
rect 16316 12004 16317 12068
rect 16251 12003 16317 12004
rect 15699 7716 15765 7717
rect 15699 7652 15700 7716
rect 15764 7652 15765 7716
rect 15699 7651 15765 7652
rect 13675 7172 13741 7173
rect 13675 7108 13676 7172
rect 13740 7108 13741 7172
rect 13675 7107 13741 7108
rect 13491 6628 13557 6629
rect 13491 6564 13492 6628
rect 13556 6564 13557 6628
rect 13491 6563 13557 6564
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 16622 5677 16682 25467
rect 24899 25260 24965 25261
rect 24899 25196 24900 25260
rect 24964 25196 24965 25260
rect 24899 25195 24965 25196
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 19931 23628 19997 23629
rect 19931 23564 19932 23628
rect 19996 23564 19997 23628
rect 19931 23563 19997 23564
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 19563 22268 19629 22269
rect 19563 22204 19564 22268
rect 19628 22204 19629 22268
rect 19563 22203 19629 22204
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 18643 20636 18709 20637
rect 18643 20572 18644 20636
rect 18708 20572 18709 20636
rect 18643 20571 18709 20572
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17171 19412 17237 19413
rect 17171 19348 17172 19412
rect 17236 19348 17237 19412
rect 17171 19347 17237 19348
rect 17174 6493 17234 19347
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18459 18052 18525 18053
rect 18459 17988 18460 18052
rect 18524 17988 18525 18052
rect 18459 17987 18525 17988
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 18462 11253 18522 17987
rect 18646 13429 18706 20571
rect 19379 20500 19445 20501
rect 19379 20436 19380 20500
rect 19444 20436 19445 20500
rect 19379 20435 19445 20436
rect 19382 15877 19442 20435
rect 19379 15876 19445 15877
rect 19379 15812 19380 15876
rect 19444 15812 19445 15876
rect 19379 15811 19445 15812
rect 18643 13428 18709 13429
rect 18643 13364 18644 13428
rect 18708 13364 18709 13428
rect 18643 13363 18709 13364
rect 19566 12885 19626 22203
rect 19747 21180 19813 21181
rect 19747 21116 19748 21180
rect 19812 21116 19813 21180
rect 19747 21115 19813 21116
rect 19750 13429 19810 21115
rect 19747 13428 19813 13429
rect 19747 13364 19748 13428
rect 19812 13364 19813 13428
rect 19747 13363 19813 13364
rect 19934 13157 19994 23563
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 24715 22676 24781 22677
rect 24715 22612 24716 22676
rect 24780 22612 24781 22676
rect 24715 22611 24781 22612
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22691 20772 22757 20773
rect 22691 20708 22692 20772
rect 22756 20708 22757 20772
rect 22691 20707 22757 20708
rect 22507 19548 22573 19549
rect 22507 19484 22508 19548
rect 22572 19484 22573 19548
rect 22507 19483 22573 19484
rect 19931 13156 19997 13157
rect 19931 13092 19932 13156
rect 19996 13092 19997 13156
rect 19931 13091 19997 13092
rect 19563 12884 19629 12885
rect 19563 12820 19564 12884
rect 19628 12820 19629 12884
rect 19563 12819 19629 12820
rect 18459 11252 18525 11253
rect 18459 11188 18460 11252
rect 18524 11188 18525 11252
rect 18459 11187 18525 11188
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 22510 7037 22570 19483
rect 22507 7036 22573 7037
rect 22507 6972 22508 7036
rect 22572 6972 22573 7036
rect 22507 6971 22573 6972
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17171 6492 17237 6493
rect 17171 6428 17172 6492
rect 17236 6428 17237 6492
rect 17171 6427 17237 6428
rect 16619 5676 16685 5677
rect 16619 5612 16620 5676
rect 16684 5612 16685 5676
rect 16619 5611 16685 5612
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 5472 18264 6496
rect 22694 5813 22754 20707
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 24718 6357 24778 22611
rect 24902 19005 24962 25195
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 24899 19004 24965 19005
rect 24899 18940 24900 19004
rect 24964 18940 24965 19004
rect 24899 18939 24965 18940
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 24715 6356 24781 6357
rect 24715 6292 24716 6356
rect 24780 6292 24781 6356
rect 24715 6291 24781 6292
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22691 5812 22757 5813
rect 22691 5748 22692 5812
rect 22756 5748 22757 5812
rect 22691 5747 22757 5748
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 33366 21725 33426 26011
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 33363 21724 33429 21725
rect 33363 21660 33364 21724
rect 33428 21660 33429 21724
rect 33363 21659 33429 21660
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1679235063
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1679235063
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1679235063
transform 1 0 5888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1679235063
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1679235063
transform 1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1679235063
transform 1 0 11776 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 10856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform 1 0 3956 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 6532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1679235063
transform 1 0 4140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1679235063
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 21068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 11960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2024 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1679235063
transform 1 0 2116 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1679235063
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 3128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1679235063
transform 1 0 2576 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _132_
timestamp 1679235063
transform 1 0 9108 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _133_
timestamp 1679235063
transform 1 0 8280 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _134_
timestamp 1679235063
transform 1 0 3312 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _135_
timestamp 1679235063
transform 1 0 5888 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_
timestamp 1679235063
transform 1 0 7636 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 36340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _139_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 38916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 37444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 35604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 36340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 38732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 33580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 34500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1679235063
transform 1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _149_
timestamp 1679235063
transform 1 0 29348 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 34868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 31464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1679235063
transform 1 0 39928 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1679235063
transform 1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _154_
timestamp 1679235063
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _155_
timestamp 1679235063
transform 1 0 33488 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 11592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 2668 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 7636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 6440 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 35788 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 26220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 4508 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 28612 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1679235063
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1679235063
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1679235063
transform 1 0 3864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 2760 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1679235063
transform 1 0 3864 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1679235063
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform 1 0 2208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1679235063
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1679235063
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1679235063
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 35420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 37628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1679235063
transform 1 0 35788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 35972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 40112 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 34868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1679235063
transform 1 0 34868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1679235063
transform 1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1679235063
transform 1 0 33948 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 36892 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 11316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10948 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1679235063
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3864 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 4048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 9292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 10856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
timestamp 1679235063
transform 1 0 22724 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 28612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
timestamp 1679235063
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 9384 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 19320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 21896 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 22080 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1679235063
transform 1 0 39284 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 36156 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold33_A
timestamp 1679235063
transform 1 0 32936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold34_A
timestamp 1679235063
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold46_A
timestamp 1679235063
transform 1 0 33212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold58_A
timestamp 1679235063
transform 1 0 36340 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold72_A
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold77_A
timestamp 1679235063
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold80_A
timestamp 1679235063
transform 1 0 40480 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold81_A
timestamp 1679235063
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold87_A
timestamp 1679235063
transform 1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold88_A
timestamp 1679235063
transform 1 0 33120 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 49128 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 4600 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 2944 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 2852 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 1472 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 4140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 34040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 37260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 39284 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 39468 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 39928 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 40480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 37812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 41124 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 38180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 42780 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 42412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 2024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 37996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 33396 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 40664 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 42964 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 49036 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 43148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 44804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1679235063
transform 1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1679235063
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1679235063
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1679235063
transform 1 0 10212 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1679235063
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1679235063
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1679235063
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1679235063
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1679235063
transform 1 0 5796 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1679235063
transform 1 0 11592 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1679235063
transform 1 0 4048 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1679235063
transform 1 0 9016 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1679235063
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 1679235063
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1679235063
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11592 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 27324 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 33580 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 27140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 33212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 33764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 31556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31740 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 30728 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29164 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 40296 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 27324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23092 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21896 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 19688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19872 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16928 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 5704 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14168 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 28520 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 35052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 5888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A1
timestamp 1679235063
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 35604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 33212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 5612 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 8280 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3864 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 14168 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 33856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 32016 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 31096 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 30912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 26588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23184 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23276 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22908 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 27876 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24472 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21344 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21160 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 29532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16744 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 37996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 10212 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 6440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 4600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 10580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 37076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 33580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 35236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8372 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4232 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4968 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5520 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5336 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 7360 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8096 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 7912 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4876 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__182 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9844 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 4140 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 9200 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 6624 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 5612 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__183
timestamp 1679235063
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 4416 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 5152 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__184
timestamp 1679235063
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 6900 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 4324 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10948 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 15272 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__185
timestamp 1679235063
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10120 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 29440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18492 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8832 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 27140 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 20884 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 25760 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 23000 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 15732 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24748 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 27600 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 14352 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17296 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9568 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 15364 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 14812 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 8740 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 13892 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 13892 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 19504 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 19504 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 25116 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 23092 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22
timestamp 1679235063
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1679235063
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1679235063
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1679235063
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1679235063
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1679235063
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1679235063
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1679235063
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1679235063
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1679235063
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1679235063
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1679235063
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1679235063
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1679235063
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1679235063
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1679235063
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1679235063
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1679235063
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1679235063
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1679235063
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_355
timestamp 1679235063
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1679235063
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1679235063
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1679235063
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1679235063
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1679235063
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1679235063
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1679235063
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1679235063
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1679235063
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1679235063
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1679235063
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1679235063
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1679235063
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1679235063
transform 1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_37
timestamp 1679235063
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1679235063
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_81
timestamp 1679235063
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1679235063
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1679235063
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1679235063
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1679235063
transform 1 0 12420 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_128
timestamp 1679235063
transform 1 0 12880 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_144
timestamp 1679235063
transform 1 0 14352 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_156
timestamp 1679235063
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1679235063
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1679235063
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_210
timestamp 1679235063
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1679235063
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1679235063
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1679235063
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1679235063
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1679235063
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1679235063
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1679235063
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1679235063
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1679235063
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1679235063
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1679235063
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1679235063
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1679235063
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1679235063
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1679235063
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1679235063
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1679235063
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1679235063
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1679235063
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1679235063
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1679235063
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1679235063
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1679235063
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1679235063
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_34
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_40
timestamp 1679235063
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1679235063
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1679235063
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp 1679235063
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_117
timestamp 1679235063
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1679235063
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1679235063
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1679235063
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1679235063
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1679235063
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1679235063
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1679235063
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1679235063
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1679235063
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1679235063
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1679235063
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1679235063
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1679235063
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1679235063
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1679235063
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1679235063
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1679235063
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1679235063
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1679235063
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1679235063
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1679235063
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1679235063
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1679235063
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_192
timestamp 1679235063
transform 1 0 18768 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_204
timestamp 1679235063
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1679235063
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1679235063
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1679235063
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1679235063
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1679235063
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1679235063
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1679235063
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1679235063
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1679235063
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1679235063
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1679235063
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1679235063
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1679235063
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1679235063
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1679235063
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1679235063
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1679235063
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1679235063
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_34
timestamp 1679235063
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_42
timestamp 1679235063
transform 1 0 4968 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_54
timestamp 1679235063
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_66
timestamp 1679235063
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1679235063
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_151
timestamp 1679235063
transform 1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_180
timestamp 1679235063
transform 1 0 17664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1679235063
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1679235063
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_210
timestamp 1679235063
transform 1 0 20424 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_222
timestamp 1679235063
transform 1 0 21528 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_234
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_240
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_258
timestamp 1679235063
transform 1 0 24840 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_270
timestamp 1679235063
transform 1 0 25944 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1679235063
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1679235063
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1679235063
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1679235063
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1679235063
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1679235063
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1679235063
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1679235063
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1679235063
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1679235063
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_22
timestamp 1679235063
transform 1 0 3128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1679235063
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1679235063
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1679235063
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_205
timestamp 1679235063
transform 1 0 19964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1679235063
transform 1 0 20700 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_227
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_233
timestamp 1679235063
transform 1 0 22540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_245
timestamp 1679235063
transform 1 0 23644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1679235063
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_304
timestamp 1679235063
transform 1 0 29072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1679235063
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1679235063
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1679235063
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1679235063
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1679235063
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1679235063
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1679235063
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1679235063
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1679235063
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1679235063
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1679235063
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1679235063
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1679235063
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1679235063
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1679235063
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1679235063
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_22
timestamp 1679235063
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1679235063
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1679235063
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_52
timestamp 1679235063
transform 1 0 5888 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_64
timestamp 1679235063
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1679235063
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1679235063
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_94
timestamp 1679235063
transform 1 0 9752 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp 1679235063
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_114
timestamp 1679235063
transform 1 0 11592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_118
timestamp 1679235063
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1679235063
transform 1 0 12696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1679235063
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1679235063
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_169
timestamp 1679235063
transform 1 0 16652 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1679235063
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_199
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_211
timestamp 1679235063
transform 1 0 20516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_223
timestamp 1679235063
transform 1 0 21620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_229
timestamp 1679235063
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_233
timestamp 1679235063
transform 1 0 22540 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_237
timestamp 1679235063
transform 1 0 22908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1679235063
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1679235063
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1679235063
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1679235063
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1679235063
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1679235063
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1679235063
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1679235063
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1679235063
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1679235063
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1679235063
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1679235063
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1679235063
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1679235063
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1679235063
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1679235063
transform 1 0 5520 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_65
timestamp 1679235063
transform 1 0 7084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_77
timestamp 1679235063
transform 1 0 8188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1679235063
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1679235063
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1679235063
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1679235063
transform 1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1679235063
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1679235063
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1679235063
transform 1 0 12788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_136
timestamp 1679235063
transform 1 0 13616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_142
timestamp 1679235063
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_146
timestamp 1679235063
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1679235063
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1679235063
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1679235063
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1679235063
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_237
timestamp 1679235063
transform 1 0 22908 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1679235063
transform 1 0 23644 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1679235063
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1679235063
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1679235063
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1679235063
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1679235063
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1679235063
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1679235063
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1679235063
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1679235063
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1679235063
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1679235063
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1679235063
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1679235063
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1679235063
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1679235063
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1679235063
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1679235063
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1679235063
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1679235063
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1679235063
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1679235063
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1679235063
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_37
timestamp 1679235063
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1679235063
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_47
timestamp 1679235063
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1679235063
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1679235063
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1679235063
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1679235063
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_103
timestamp 1679235063
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1679235063
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1679235063
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1679235063
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1679235063
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1679235063
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1679235063
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1679235063
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1679235063
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1679235063
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1679235063
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1679235063
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1679235063
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1679235063
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1679235063
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1679235063
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1679235063
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1679235063
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1679235063
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp 1679235063
transform 1 0 3036 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1679235063
transform 1 0 4232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp 1679235063
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1679235063
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1679235063
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 1679235063
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_73
timestamp 1679235063
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1679235063
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_88
timestamp 1679235063
transform 1 0 9200 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1679235063
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1679235063
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1679235063
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1679235063
transform 1 0 13800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1679235063
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1679235063
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1679235063
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_174
timestamp 1679235063
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_186
timestamp 1679235063
transform 1 0 18216 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_198
timestamp 1679235063
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_210
timestamp 1679235063
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp 1679235063
transform 1 0 22172 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_250
timestamp 1679235063
transform 1 0 24104 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_254
timestamp 1679235063
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_266
timestamp 1679235063
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1679235063
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1679235063
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1679235063
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1679235063
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1679235063
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1679235063
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1679235063
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1679235063
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1679235063
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1679235063
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1679235063
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1679235063
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1679235063
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1679235063
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1679235063
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1679235063
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1679235063
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1679235063
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1679235063
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1679235063
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1679235063
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_8
timestamp 1679235063
transform 1 0 1840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1679235063
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1679235063
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1679235063
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1679235063
transform 1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1679235063
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1679235063
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_69
timestamp 1679235063
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1679235063
transform 1 0 7820 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_91
timestamp 1679235063
transform 1 0 9476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1679235063
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1679235063
transform 1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1679235063
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1679235063
transform 1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1679235063
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_152
timestamp 1679235063
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1679235063
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1679235063
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_178
timestamp 1679235063
transform 1 0 17480 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_184
timestamp 1679235063
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1679235063
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1679235063
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1679235063
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1679235063
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1679235063
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1679235063
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1679235063
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1679235063
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1679235063
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1679235063
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1679235063
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1679235063
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1679235063
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1679235063
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1679235063
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1679235063
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1679235063
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1679235063
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1679235063
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1679235063
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1679235063
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1679235063
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1679235063
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1679235063
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1679235063
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_8
timestamp 1679235063
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1679235063
transform 1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1679235063
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1679235063
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1679235063
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1679235063
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1679235063
transform 1 0 10672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1679235063
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1679235063
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1679235063
transform 1 0 14260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1679235063
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1679235063
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_171
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1679235063
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp 1679235063
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_198
timestamp 1679235063
transform 1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_202
timestamp 1679235063
transform 1 0 19688 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1679235063
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1679235063
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1679235063
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1679235063
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1679235063
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1679235063
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1679235063
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1679235063
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1679235063
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1679235063
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1679235063
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1679235063
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1679235063
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1679235063
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1679235063
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1679235063
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1679235063
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1679235063
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1679235063
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1679235063
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1679235063
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1679235063
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1679235063
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1679235063
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1679235063
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_8
timestamp 1679235063
transform 1 0 1840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_14
timestamp 1679235063
transform 1 0 2392 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_35
timestamp 1679235063
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1679235063
transform 1 0 4784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1679235063
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1679235063
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1679235063
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1679235063
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_97
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1679235063
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1679235063
transform 1 0 12420 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1679235063
transform 1 0 12788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1679235063
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1679235063
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1679235063
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_206
timestamp 1679235063
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_217
timestamp 1679235063
transform 1 0 21068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_229
timestamp 1679235063
transform 1 0 22172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_241
timestamp 1679235063
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1679235063
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1679235063
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_277
timestamp 1679235063
transform 1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_285
timestamp 1679235063
transform 1 0 27324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_295
timestamp 1679235063
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1679235063
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1679235063
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1679235063
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1679235063
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1679235063
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1679235063
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1679235063
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1679235063
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1679235063
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1679235063
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1679235063
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1679235063
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1679235063
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1679235063
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1679235063
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1679235063
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1679235063
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1679235063
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1679235063
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1679235063
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1679235063
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1679235063
transform 1 0 3036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1679235063
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1679235063
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_63
timestamp 1679235063
transform 1 0 6900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1679235063
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1679235063
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1679235063
transform 1 0 14076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1679235063
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1679235063
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_204
timestamp 1679235063
transform 1 0 19872 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_216
timestamp 1679235063
transform 1 0 20976 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_235
timestamp 1679235063
transform 1 0 22724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_247
timestamp 1679235063
transform 1 0 23828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_259
timestamp 1679235063
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1679235063
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1679235063
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_291
timestamp 1679235063
transform 1 0 27876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_303
timestamp 1679235063
transform 1 0 28980 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_315
timestamp 1679235063
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp 1679235063
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1679235063
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1679235063
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1679235063
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1679235063
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1679235063
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1679235063
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1679235063
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1679235063
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1679235063
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1679235063
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1679235063
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1679235063
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1679235063
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1679235063
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1679235063
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1679235063
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_23
timestamp 1679235063
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_35
timestamp 1679235063
transform 1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1679235063
transform 1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1679235063
transform 1 0 5428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_56
timestamp 1679235063
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1679235063
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1679235063
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1679235063
transform 1 0 11316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1679235063
transform 1 0 13248 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1679235063
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_171
timestamp 1679235063
transform 1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_220
timestamp 1679235063
transform 1 0 21344 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1679235063
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1679235063
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1679235063
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1679235063
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1679235063
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1679235063
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1679235063
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1679235063
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1679235063
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1679235063
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1679235063
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1679235063
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1679235063
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1679235063
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1679235063
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1679235063
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1679235063
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1679235063
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1679235063
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1679235063
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1679235063
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1679235063
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1679235063
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1679235063
transform 1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_14
timestamp 1679235063
transform 1 0 2392 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_26
timestamp 1679235063
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1679235063
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1679235063
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1679235063
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1679235063
transform 1 0 9844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1679235063
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1679235063
transform 1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1679235063
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1679235063
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_227
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1679235063
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1679235063
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1679235063
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1679235063
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1679235063
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1679235063
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1679235063
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1679235063
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1679235063
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1679235063
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1679235063
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1679235063
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1679235063
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1679235063
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1679235063
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1679235063
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1679235063
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1679235063
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1679235063
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1679235063
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1679235063
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1679235063
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1679235063
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1679235063
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1679235063
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1679235063
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_20
timestamp 1679235063
transform 1 0 2944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_35
timestamp 1679235063
transform 1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_40
timestamp 1679235063
transform 1 0 4784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1679235063
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1679235063
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1679235063
transform 1 0 11224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1679235063
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1679235063
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_169
timestamp 1679235063
transform 1 0 16652 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_173
timestamp 1679235063
transform 1 0 17020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_211
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_235
timestamp 1679235063
transform 1 0 22724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_247
timestamp 1679235063
transform 1 0 23828 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1679235063
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1679235063
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1679235063
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1679235063
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1679235063
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1679235063
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1679235063
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1679235063
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1679235063
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1679235063
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1679235063
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1679235063
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1679235063
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1679235063
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1679235063
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1679235063
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1679235063
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1679235063
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1679235063
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1679235063
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1679235063
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1679235063
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1679235063
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_14
timestamp 1679235063
transform 1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1679235063
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1679235063
transform 1 0 3772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1679235063
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_63
timestamp 1679235063
transform 1 0 6900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_67
timestamp 1679235063
transform 1 0 7268 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1679235063
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1679235063
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1679235063
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_173
timestamp 1679235063
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1679235063
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1679235063
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_257
timestamp 1679235063
transform 1 0 24748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1679235063
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1679235063
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1679235063
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1679235063
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1679235063
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1679235063
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1679235063
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1679235063
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1679235063
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1679235063
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1679235063
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1679235063
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1679235063
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1679235063
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1679235063
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1679235063
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1679235063
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1679235063
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1679235063
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1679235063
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1679235063
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1679235063
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1679235063
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1679235063
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_34
timestamp 1679235063
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1679235063
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1679235063
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1679235063
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_102
timestamp 1679235063
transform 1 0 10488 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1679235063
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1679235063
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1679235063
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1679235063
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1679235063
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_203
timestamp 1679235063
transform 1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_264
timestamp 1679235063
transform 1 0 25392 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1679235063
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1679235063
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1679235063
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1679235063
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1679235063
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1679235063
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1679235063
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1679235063
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1679235063
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1679235063
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1679235063
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1679235063
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1679235063
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1679235063
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1679235063
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1679235063
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1679235063
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1679235063
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1679235063
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1679235063
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1679235063
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1679235063
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1679235063
transform 1 0 3864 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1679235063
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_61
timestamp 1679235063
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_72
timestamp 1679235063
transform 1 0 7728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1679235063
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1679235063
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_115
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_118
timestamp 1679235063
transform 1 0 11960 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_121
timestamp 1679235063
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1679235063
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1679235063
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_171
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_183
timestamp 1679235063
transform 1 0 17940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1679235063
transform 1 0 19136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_211
timestamp 1679235063
transform 1 0 20516 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_218
timestamp 1679235063
transform 1 0 21160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1679235063
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1679235063
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1679235063
transform 1 0 24840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1679235063
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1679235063
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1679235063
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1679235063
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1679235063
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1679235063
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1679235063
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1679235063
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1679235063
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1679235063
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1679235063
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1679235063
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1679235063
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1679235063
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1679235063
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1679235063
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1679235063
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1679235063
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1679235063
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1679235063
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1679235063
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1679235063
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_34
timestamp 1679235063
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1679235063
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1679235063
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1679235063
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1679235063
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_115
timestamp 1679235063
transform 1 0 11684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1679235063
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_202
timestamp 1679235063
transform 1 0 19688 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1679235063
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1679235063
transform 1 0 22080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_235
timestamp 1679235063
transform 1 0 22724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_239
timestamp 1679235063
transform 1 0 23092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1679235063
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_276
timestamp 1679235063
transform 1 0 26496 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_288
timestamp 1679235063
transform 1 0 27600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1679235063
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1679235063
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1679235063
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1679235063
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1679235063
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1679235063
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1679235063
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1679235063
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1679235063
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1679235063
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1679235063
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1679235063
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1679235063
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1679235063
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1679235063
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1679235063
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1679235063
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1679235063
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1679235063
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1679235063
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1679235063
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1679235063
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_125
timestamp 1679235063
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1679235063
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_150
timestamp 1679235063
transform 1 0 14904 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_154
timestamp 1679235063
transform 1 0 15272 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_164
timestamp 1679235063
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1679235063
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1679235063
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_216
timestamp 1679235063
transform 1 0 20976 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1679235063
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1679235063
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1679235063
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1679235063
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1679235063
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1679235063
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1679235063
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1679235063
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1679235063
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1679235063
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1679235063
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1679235063
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1679235063
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1679235063
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1679235063
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1679235063
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1679235063
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1679235063
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1679235063
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1679235063
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1679235063
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1679235063
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1679235063
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_31
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1679235063
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1679235063
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1679235063
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1679235063
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_144
timestamp 1679235063
transform 1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_191
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1679235063
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_225
timestamp 1679235063
transform 1 0 21804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1679235063
transform 1 0 22080 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1679235063
transform 1 0 24932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_272
timestamp 1679235063
transform 1 0 26128 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_284
timestamp 1679235063
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_296
timestamp 1679235063
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1679235063
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1679235063
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1679235063
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1679235063
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1679235063
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1679235063
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1679235063
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1679235063
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1679235063
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1679235063
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1679235063
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1679235063
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1679235063
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1679235063
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1679235063
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1679235063
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1679235063
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_25
timestamp 1679235063
transform 1 0 3404 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1679235063
transform 1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1679235063
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1679235063
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1679235063
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1679235063
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_119
timestamp 1679235063
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1679235063
transform 1 0 13248 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_136
timestamp 1679235063
transform 1 0 13616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_174
timestamp 1679235063
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1679235063
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_235
timestamp 1679235063
transform 1 0 22724 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_250
timestamp 1679235063
transform 1 0 24104 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1679235063
transform 1 0 24656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1679235063
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1679235063
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1679235063
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1679235063
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1679235063
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1679235063
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1679235063
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1679235063
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1679235063
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1679235063
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1679235063
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1679235063
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1679235063
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1679235063
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1679235063
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1679235063
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1679235063
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1679235063
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1679235063
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1679235063
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1679235063
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1679235063
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1679235063
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1679235063
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1679235063
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_66
timestamp 1679235063
transform 1 0 7176 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1679235063
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1679235063
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1679235063
transform 1 0 10488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1679235063
transform 1 0 10856 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_116
timestamp 1679235063
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1679235063
transform 1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1679235063
transform 1 0 13340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1679235063
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1679235063
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1679235063
transform 1 0 16744 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_199
timestamp 1679235063
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_211
timestamp 1679235063
transform 1 0 20516 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1679235063
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_237
timestamp 1679235063
transform 1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1679235063
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1679235063
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1679235063
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_296
timestamp 1679235063
transform 1 0 28336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1679235063
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1679235063
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1679235063
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1679235063
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1679235063
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1679235063
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1679235063
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1679235063
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1679235063
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1679235063
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1679235063
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1679235063
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1679235063
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1679235063
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1679235063
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1679235063
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1679235063
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1679235063
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1679235063
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1679235063
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1679235063
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1679235063
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_89
timestamp 1679235063
transform 1 0 9292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_96
timestamp 1679235063
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_107
timestamp 1679235063
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1679235063
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1679235063
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_186
timestamp 1679235063
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_192
timestamp 1679235063
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_202
timestamp 1679235063
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1679235063
transform 1 0 20884 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1679235063
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_243
timestamp 1679235063
transform 1 0 23460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1679235063
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_291
timestamp 1679235063
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_303
timestamp 1679235063
transform 1 0 28980 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_311
timestamp 1679235063
transform 1 0 29716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_323
timestamp 1679235063
transform 1 0 30820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1679235063
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1679235063
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1679235063
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1679235063
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1679235063
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1679235063
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1679235063
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1679235063
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1679235063
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1679235063
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1679235063
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1679235063
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1679235063
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1679235063
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1679235063
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1679235063
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1679235063
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1679235063
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_51
timestamp 1679235063
transform 1 0 5796 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_56
timestamp 1679235063
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1679235063
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1679235063
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1679235063
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1679235063
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1679235063
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_166
timestamp 1679235063
transform 1 0 16376 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1679235063
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_189
timestamp 1679235063
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1679235063
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_235
timestamp 1679235063
transform 1 0 22724 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_239
timestamp 1679235063
transform 1 0 23092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_266
timestamp 1679235063
transform 1 0 25576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1679235063
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1679235063
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1679235063
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1679235063
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1679235063
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1679235063
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1679235063
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1679235063
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1679235063
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1679235063
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1679235063
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1679235063
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1679235063
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1679235063
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1679235063
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1679235063
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1679235063
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1679235063
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1679235063
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1679235063
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1679235063
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1679235063
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_60
timestamp 1679235063
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_119
timestamp 1679235063
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1679235063
transform 1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_140
timestamp 1679235063
transform 1 0 13984 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1679235063
transform 1 0 18032 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1679235063
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_209
timestamp 1679235063
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1679235063
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_227
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_238
timestamp 1679235063
transform 1 0 23000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_242
timestamp 1679235063
transform 1 0 23368 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1679235063
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1679235063
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1679235063
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_311
timestamp 1679235063
transform 1 0 29716 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_315
timestamp 1679235063
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_327
timestamp 1679235063
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1679235063
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1679235063
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1679235063
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1679235063
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1679235063
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1679235063
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1679235063
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1679235063
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1679235063
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1679235063
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1679235063
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1679235063
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1679235063
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1679235063
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1679235063
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1679235063
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1679235063
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1679235063
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_80
timestamp 1679235063
transform 1 0 8464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1679235063
transform 1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_135
timestamp 1679235063
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1679235063
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1679235063
transform 1 0 14996 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1679235063
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1679235063
transform 1 0 18124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1679235063
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_199
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1679235063
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 1679235063
transform 1 0 21528 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_257
timestamp 1679235063
transform 1 0 24748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1679235063
transform 1 0 26772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_303
timestamp 1679235063
transform 1 0 28980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1679235063
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_320
timestamp 1679235063
transform 1 0 30544 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_330
timestamp 1679235063
transform 1 0 31464 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_342
timestamp 1679235063
transform 1 0 32568 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_354
timestamp 1679235063
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1679235063
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1679235063
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1679235063
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1679235063
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1679235063
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1679235063
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1679235063
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1679235063
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1679235063
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1679235063
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1679235063
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1679235063
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1679235063
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1679235063
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1679235063
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_79
timestamp 1679235063
transform 1 0 8372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1679235063
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_107
timestamp 1679235063
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_122
timestamp 1679235063
transform 1 0 12328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1679235063
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_150
timestamp 1679235063
transform 1 0 14904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_163
timestamp 1679235063
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_194
timestamp 1679235063
transform 1 0 18952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1679235063
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_212
timestamp 1679235063
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1679235063
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_274
timestamp 1679235063
transform 1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1679235063
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_286
timestamp 1679235063
transform 1 0 27416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_290
timestamp 1679235063
transform 1 0 27784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1679235063
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_326
timestamp 1679235063
transform 1 0 31096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1679235063
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_339
timestamp 1679235063
transform 1 0 32292 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_351
timestamp 1679235063
transform 1 0 33396 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_363
timestamp 1679235063
transform 1 0 34500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_375
timestamp 1679235063
transform 1 0 35604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1679235063
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1679235063
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1679235063
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1679235063
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1679235063
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1679235063
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1679235063
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1679235063
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1679235063
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1679235063
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1679235063
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1679235063
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1679235063
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1679235063
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_33
timestamp 1679235063
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_44
timestamp 1679235063
transform 1 0 5152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_68
timestamp 1679235063
transform 1 0 7360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1679235063
transform 1 0 10028 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_112
timestamp 1679235063
transform 1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_129
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1679235063
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1679235063
transform 1 0 14812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_173
timestamp 1679235063
transform 1 0 17020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1679235063
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1679235063
transform 1 0 20608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1679235063
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1679235063
transform 1 0 24840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1679235063
transform 1 0 25208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_284
timestamp 1679235063
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1679235063
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_304
timestamp 1679235063
transform 1 0 29072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1679235063
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_332
timestamp 1679235063
transform 1 0 31648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_338
timestamp 1679235063
transform 1 0 32200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_344
timestamp 1679235063
transform 1 0 32752 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1679235063
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1679235063
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1679235063
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1679235063
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1679235063
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1679235063
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1679235063
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1679235063
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1679235063
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1679235063
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1679235063
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1679235063
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1679235063
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1679235063
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1679235063
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_30
timestamp 1679235063
transform 1 0 3864 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_63
timestamp 1679235063
transform 1 0 6900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_87
timestamp 1679235063
transform 1 0 9108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1679235063
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 1679235063
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1679235063
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_163
timestamp 1679235063
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_175
timestamp 1679235063
transform 1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1679235063
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_198
timestamp 1679235063
transform 1 0 19320 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_230
timestamp 1679235063
transform 1 0 22264 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1679235063
transform 1 0 24472 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1679235063
transform 1 0 24840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_270
timestamp 1679235063
transform 1 0 25944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1679235063
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_292
timestamp 1679235063
transform 1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1679235063
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_328
timestamp 1679235063
transform 1 0 31280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_343
timestamp 1679235063
transform 1 0 32660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_351
timestamp 1679235063
transform 1 0 33396 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_355
timestamp 1679235063
transform 1 0 33764 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_367
timestamp 1679235063
transform 1 0 34868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_379
timestamp 1679235063
transform 1 0 35972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1679235063
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1679235063
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1679235063
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1679235063
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1679235063
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1679235063
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1679235063
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1679235063
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1679235063
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1679235063
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1679235063
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1679235063
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1679235063
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_36
timestamp 1679235063
transform 1 0 4416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_40
timestamp 1679235063
transform 1 0 4784 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1679235063
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1679235063
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1679235063
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1679235063
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1679235063
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1679235063
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1679235063
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 1679235063
transform 1 0 16928 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1679235063
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_203
timestamp 1679235063
transform 1 0 19780 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1679235063
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_234
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_247
timestamp 1679235063
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1679235063
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1679235063
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1679235063
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 1679235063
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_334
timestamp 1679235063
transform 1 0 31832 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_346
timestamp 1679235063
transform 1 0 32936 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_350
timestamp 1679235063
transform 1 0 33304 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1679235063
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_369
timestamp 1679235063
transform 1 0 35052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_381
timestamp 1679235063
transform 1 0 36156 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_393
timestamp 1679235063
transform 1 0 37260 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_405
timestamp 1679235063
transform 1 0 38364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_417
timestamp 1679235063
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1679235063
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1679235063
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1679235063
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1679235063
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1679235063
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1679235063
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1679235063
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1679235063
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1679235063
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1679235063
transform 1 0 8372 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_101
timestamp 1679235063
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_105
timestamp 1679235063
transform 1 0 10764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1679235063
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_133
timestamp 1679235063
transform 1 0 13340 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1679235063
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1679235063
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_182
timestamp 1679235063
transform 1 0 17848 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1679235063
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_235
timestamp 1679235063
transform 1 0 22724 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_248
timestamp 1679235063
transform 1 0 23920 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_272
timestamp 1679235063
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1679235063
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_296
timestamp 1679235063
transform 1 0 28336 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1679235063
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1679235063
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_347
timestamp 1679235063
transform 1 0 33028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_351
timestamp 1679235063
transform 1 0 33396 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1679235063
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_365
timestamp 1679235063
transform 1 0 34684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_381
timestamp 1679235063
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1679235063
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1679235063
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1679235063
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1679235063
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1679235063
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1679235063
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1679235063
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1679235063
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1679235063
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1679235063
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1679235063
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1679235063
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_54
timestamp 1679235063
transform 1 0 6072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1679235063
transform 1 0 8096 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1679235063
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_111
timestamp 1679235063
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp 1679235063
transform 1 0 11776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_146
timestamp 1679235063
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_157
timestamp 1679235063
transform 1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1679235063
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_190
timestamp 1679235063
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_247
timestamp 1679235063
transform 1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1679235063
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1679235063
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_302
timestamp 1679235063
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_319
timestamp 1679235063
transform 1 0 30452 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_331
timestamp 1679235063
transform 1 0 31556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_335
timestamp 1679235063
transform 1 0 31924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_341
timestamp 1679235063
transform 1 0 32476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_355
timestamp 1679235063
transform 1 0 33764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1679235063
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_371
timestamp 1679235063
transform 1 0 35236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_379
timestamp 1679235063
transform 1 0 35972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1679235063
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_395
timestamp 1679235063
transform 1 0 37444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_407
timestamp 1679235063
transform 1 0 38548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1679235063
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1679235063
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1679235063
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1679235063
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1679235063
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1679235063
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1679235063
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1679235063
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1679235063
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_71
timestamp 1679235063
transform 1 0 7636 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_94
timestamp 1679235063
transform 1 0 9752 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1679235063
transform 1 0 10212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_116
timestamp 1679235063
transform 1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_127
timestamp 1679235063
transform 1 0 12788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_151
timestamp 1679235063
transform 1 0 14996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1679235063
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1679235063
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1679235063
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1679235063
transform 1 0 20424 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1679235063
transform 1 0 26404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1679235063
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1679235063
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1679235063
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1679235063
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_347
timestamp 1679235063
transform 1 0 33028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_354
timestamp 1679235063
transform 1 0 33672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_360
timestamp 1679235063
transform 1 0 34224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1679235063
transform 1 0 34868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_382
timestamp 1679235063
transform 1 0 36248 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1679235063
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_407
timestamp 1679235063
transform 1 0 38548 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_419
timestamp 1679235063
transform 1 0 39652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_431
timestamp 1679235063
transform 1 0 40756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_443
timestamp 1679235063
transform 1 0 41860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1679235063
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1679235063
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1679235063
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1679235063
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1679235063
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1679235063
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1679235063
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1679235063
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1679235063
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1679235063
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1679235063
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1679235063
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1679235063
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_225
timestamp 1679235063
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1679235063
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1679235063
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_300
timestamp 1679235063
transform 1 0 28704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_311
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_323
timestamp 1679235063
transform 1 0 30820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_335
timestamp 1679235063
transform 1 0 31924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_347
timestamp 1679235063
transform 1 0 33028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_359
timestamp 1679235063
transform 1 0 34132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1679235063
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_371
timestamp 1679235063
transform 1 0 35236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_379
timestamp 1679235063
transform 1 0 35972 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_385
timestamp 1679235063
transform 1 0 36524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_392
timestamp 1679235063
transform 1 0 37168 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_399
timestamp 1679235063
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_406
timestamp 1679235063
transform 1 0 38456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_413
timestamp 1679235063
transform 1 0 39100 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_417
timestamp 1679235063
transform 1 0 39468 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1679235063
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1679235063
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1679235063
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1679235063
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1679235063
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1679235063
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1679235063
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1679235063
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_25
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_70
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1679235063
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_144
timestamp 1679235063
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1679235063
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1679235063
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1679235063
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_291
timestamp 1679235063
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_295
timestamp 1679235063
transform 1 0 28244 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1679235063
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_329
timestamp 1679235063
transform 1 0 31372 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1679235063
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_347
timestamp 1679235063
transform 1 0 33028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_351
timestamp 1679235063
transform 1 0 33396 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_357
timestamp 1679235063
transform 1 0 33948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_371
timestamp 1679235063
transform 1 0 35236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_379
timestamp 1679235063
transform 1 0 35972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_387
timestamp 1679235063
transform 1 0 36708 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1679235063
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_397
timestamp 1679235063
transform 1 0 37628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_420
timestamp 1679235063
transform 1 0 39744 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_430
timestamp 1679235063
transform 1 0 40664 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_434
timestamp 1679235063
transform 1 0 41032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_437
timestamp 1679235063
transform 1 0 41308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1679235063
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1679235063
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1679235063
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1679235063
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1679235063
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1679235063
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1679235063
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1679235063
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1679235063
transform 1 0 9200 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1679235063
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_135
timestamp 1679235063
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_152
timestamp 1679235063
transform 1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1679235063
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1679235063
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1679235063
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_281
timestamp 1679235063
transform 1 0 26956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_304
timestamp 1679235063
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1679235063
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_343
timestamp 1679235063
transform 1 0 32660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_355
timestamp 1679235063
transform 1 0 33764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1679235063
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_370
timestamp 1679235063
transform 1 0 35144 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_384
timestamp 1679235063
transform 1 0 36432 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_391
timestamp 1679235063
transform 1 0 37076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_399
timestamp 1679235063
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_407
timestamp 1679235063
transform 1 0 38548 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_415
timestamp 1679235063
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1679235063
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_426
timestamp 1679235063
transform 1 0 40296 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_433
timestamp 1679235063
transform 1 0 40940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_440
timestamp 1679235063
transform 1 0 41584 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_447
timestamp 1679235063
transform 1 0 42228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_451
timestamp 1679235063
transform 1 0 42596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_463
timestamp 1679235063
transform 1 0 43700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1679235063
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1679235063
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1679235063
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1679235063
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1679235063
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 1679235063
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_171
timestamp 1679235063
transform 1 0 16836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1679235063
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_213
timestamp 1679235063
transform 1 0 20700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1679235063
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1679235063
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1679235063
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1679235063
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1679235063
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_325
timestamp 1679235063
transform 1 0 31004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_332
timestamp 1679235063
transform 1 0 31648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_347
timestamp 1679235063
transform 1 0 33028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_359
timestamp 1679235063
transform 1 0 34132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_371
timestamp 1679235063
transform 1 0 35236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1679235063
transform 1 0 35972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1679235063
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1679235063
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_398
timestamp 1679235063
transform 1 0 37720 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1679235063
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_413
timestamp 1679235063
transform 1 0 39100 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_419
timestamp 1679235063
transform 1 0 39652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_426
timestamp 1679235063
transform 1 0 40296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1679235063
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_459
timestamp 1679235063
transform 1 0 43332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_465
timestamp 1679235063
transform 1 0 43884 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_473
timestamp 1679235063
transform 1 0 44620 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_477
timestamp 1679235063
transform 1 0 44988 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_487
timestamp 1679235063
transform 1 0 45908 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_495
timestamp 1679235063
transform 1 0 46644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1679235063
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_507
timestamp 1679235063
transform 1 0 47748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_515
timestamp 1679235063
transform 1 0 48484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_520
timestamp 1679235063
transform 1 0 48944 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_524
timestamp 1679235063
transform 1 0 49312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1679235063
transform 1 0 4416 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_120
timestamp 1679235063
transform 1 0 12144 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_191
timestamp 1679235063
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1679235063
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_287
timestamp 1679235063
transform 1 0 27508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_298
timestamp 1679235063
transform 1 0 28520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1679235063
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_333
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_347
timestamp 1679235063
transform 1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_359
timestamp 1679235063
transform 1 0 34132 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1679235063
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_375
timestamp 1679235063
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_383
timestamp 1679235063
transform 1 0 36340 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_390
timestamp 1679235063
transform 1 0 36984 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_399
timestamp 1679235063
transform 1 0 37812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_403
timestamp 1679235063
transform 1 0 38180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_409
timestamp 1679235063
transform 1 0 38732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_417
timestamp 1679235063
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_426
timestamp 1679235063
transform 1 0 40296 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_434
timestamp 1679235063
transform 1 0 41032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1679235063
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_471
timestamp 1679235063
transform 1 0 44436 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1679235063
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1679235063
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1679235063
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1679235063
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1679235063
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_519
timestamp 1679235063
transform 1 0 48852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_523
timestamp 1679235063
transform 1 0 49220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 33396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 27968 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 13064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold6
timestamp 1679235063
transform 1 0 11684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold9
timestamp 1679235063
transform 1 0 32292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 27600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 4416 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold12
timestamp 1679235063
transform 1 0 34316 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 2760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold14
timestamp 1679235063
transform 1 0 3496 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 14260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold16
timestamp 1679235063
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold17
timestamp 1679235063
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold18
timestamp 1679235063
transform 1 0 33396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold20
timestamp 1679235063
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 10672 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1679235063
transform 1 0 5520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold23
timestamp 1679235063
transform 1 0 32292 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold24
timestamp 1679235063
transform 1 0 33672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold25
timestamp 1679235063
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 19596 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 22172 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 30820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 28060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold30
timestamp 1679235063
transform 1 0 6808 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold31
timestamp 1679235063
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold33
timestamp 1679235063
transform 1 0 32476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold34
timestamp 1679235063
transform 1 0 1656 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold35
timestamp 1679235063
transform 1 0 30544 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 23092 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold37
timestamp 1679235063
transform 1 0 3128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1679235063
transform 1 0 27232 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1679235063
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 20240 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold41
timestamp 1679235063
transform 1 0 5612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 12788 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 17204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 12604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold46
timestamp 1679235063
transform 1 0 32844 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 20792 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 16652 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 12880 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 31004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 30912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold58
timestamp 1679235063
transform 1 0 34316 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 33028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 9292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 11500 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 15364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold65
timestamp 1679235063
transform 1 0 32292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 4232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold67
timestamp 1679235063
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 27140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 28152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1679235063
transform 1 0 6716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold72
timestamp 1679235063
transform 1 0 34132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold73
timestamp 1679235063
transform 1 0 31924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 31188 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1679235063
transform 1 0 29716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 28244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold77
timestamp 1679235063
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform 1 0 27140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1679235063
transform 1 0 32292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold80
timestamp 1679235063
transform 1 0 34868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold81
timestamp 1679235063
transform 1 0 3496 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 21712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 26496 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold86
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold87
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold88
timestamp 1679235063
transform 1 0 32200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1679235063
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 21988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform 1 0 7268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1679235063
transform 1 0 18584 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold95
timestamp 1679235063
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 23276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 25208 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 48668 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1679235063
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1679235063
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 6440 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 2852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1679235063
transform 1 0 1564 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 2852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1679235063
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1679235063
transform 1 0 3312 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1679235063
transform 1 0 35512 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1679235063
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 38088 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 36800 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1679235063
transform 1 0 35972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1679235063
transform 1 0 36340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 31372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1679235063
transform 1 0 37444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 40664 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 36616 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 41308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 38180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1679235063
transform 1 0 38364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1679235063
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 40664 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1679235063
transform 1 0 41216 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 41952 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1679235063
transform 1 0 1564 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 34132 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 34868 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1679235063
transform 1 0 36708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1679235063
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1679235063
transform 1 0 48484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1679235063
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 44252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 7084 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 5796 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 17112 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 17020 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 7912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24932 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20148 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21160 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18860 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24288 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25944 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27232 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28336 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28428 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28336 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24748 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37904 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27876 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22356 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19504 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20884 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21068 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23000 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16008 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14812 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16192 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14536 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12144 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11408 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11592 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8556 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7268 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5520 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4232 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6256 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7820 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9384 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12420 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13156 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13708 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 15180 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16284 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18124 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 31004 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 28428 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__186
timestamp 1679235063
transform 1 0 27232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__145
timestamp 1679235063
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 34316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23644 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__154
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14536 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 33396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12512 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__187
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14720 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__188
timestamp 1679235063
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__189
timestamp 1679235063
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 32292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__190
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__143
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__144
timestamp 1679235063
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22448 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__146
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27692 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__147
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30544 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  sb_8__0_.mux_left_track_35.mux_l2_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__148
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29992 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__149
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__150
timestamp 1679235063
transform 1 0 32200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 27600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__151
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22172 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 27232 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__156
timestamp 1679235063
transform 1 0 19504 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23644 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22356 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 26404 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 13064 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__162
timestamp 1679235063
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 25944 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23184 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17112 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__173
timestamp 1679235063
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23552 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__180
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14352 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19688 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24748 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14352 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__181
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 20148 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14352 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__157
timestamp 1679235063
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 22448 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__158
timestamp 1679235063
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17204 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10212 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__159
timestamp 1679235063
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29716 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__160
timestamp 1679235063
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12880 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14076 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__161
timestamp 1679235063
transform 1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15916 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14720 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14996 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__164
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15364 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__165
timestamp 1679235063
transform 1 0 7820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18400 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__166
timestamp 1679235063
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__167
timestamp 1679235063
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12144 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__168
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 26404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__169
timestamp 1679235063
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12420 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10580 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__170
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__171
timestamp 1679235063
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 8464 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6624 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__172
timestamp 1679235063
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6716 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6716 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__175
timestamp 1679235063
transform 1 0 35972 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9752 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__176
timestamp 1679235063
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 36800 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__177
timestamp 1679235063
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19780 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__178
timestamp 1679235063
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15272 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__179
timestamp 1679235063
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 34868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 18538 4828 18538 4828 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 16882 4998 16882 4998 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 15456 4658 15456 4658 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 14398 5644 14398 5644 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20838 17136 20838 17136 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 7958 7922 7958 7922 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal2 20746 15028 20746 15028 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 10718 14042 10718 14042 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal2 10902 9792 10902 9792 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 6532 10982 6532 10982 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 6164 16014 6164 16014 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 5474 14926 5474 14926 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal2 6026 13056 6026 13056 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 8326 11526 8326 11526 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal2 7682 13889 7682 13889 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal2 12558 16303 12558 16303 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 7590 12784 7590 12784 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 8188 17714 8188 17714 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 7406 17068 7406 17068 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 5704 20366 5704 20366 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal2 8602 14960 8602 14960 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9890 8738 9890 8738 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15134 6800 15134 6800 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 8418 14042 8418 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9913 15538 9913 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10258 15470 10258 15470 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12604 12614 12604 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8004 14042 8004 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9706 13226 9706 13226 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9982 8534 9982 8534 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10350 8602 10350 8602 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12144 8874 12144 8874 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4186 14756 4186 14756 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6808 10778 6808 10778 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 11914 5712 11914 5712 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 5014 18224 5014 18224 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6716 15538 6716 15538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7314 15470 7314 15470 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10258 14246 10258 14246 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 4784 13362 4784 13362 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 5152 13294 5152 13294 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6624 10234 6624 10234 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 5704 13158 5704 13158 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 4784 13430 4784 13430 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4830 15402 4830 15402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9292 9894 9292 9894 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13041 5678 13041 5678 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 5566 16218 5566 16218 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7038 13974 7038 13974 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7314 14144 7314 14144 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10212 14790 10212 14790 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7084 12818 7084 12818 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7130 12954 7130 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8280 11322 8280 11322 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14030 15062 14030 15062 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8050 10098 8050 10098 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 8280 17306 8280 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6026 18326 6026 18326 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel via3 5267 13668 5267 13668 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 6394 17306 6394 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7130 17068 7130 17068 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7728 15674 7728 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 9890 14892 9890 14892 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 6624 17034 6624 17034 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6578 16422 6578 16422 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8970 14586 8970 14586 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12374 18394 12374 18394 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 5750 19312 5750 19312 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14306 4658 14306 4658 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 17296 3094 17296 3094 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 27209 4726 27209 4726 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 20746 5882 20746 5882 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 15594 4046 15594 4046 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 25231 4794 25231 4794 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 24058 8534 24058 8534 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 13248 3094 13248 3094 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 22977 5338 22977 5338 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 14950 5610 14950 5610 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 24886 5270 24886 5270 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 2944 2414 2944 2414 0 ccff_head
rlabel metal2 48898 25007 48898 25007 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2254 22348 2254 22348 0 ccff_tail_0
rlabel metal2 3358 2176 3358 2176 0 chanx_left_in[0]
rlabel metal3 1142 5644 1142 5644 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 4232 4590 4232 4590 0 chanx_left_in[12]
rlabel metal3 2668 6800 2668 6800 0 chanx_left_in[13]
rlabel metal1 4462 5202 4462 5202 0 chanx_left_in[14]
rlabel metal1 4922 6290 4922 6290 0 chanx_left_in[15]
rlabel metal1 4554 5678 4554 5678 0 chanx_left_in[16]
rlabel metal1 3818 5202 3818 5202 0 chanx_left_in[17]
rlabel metal2 6670 7548 6670 7548 0 chanx_left_in[18]
rlabel metal2 2714 7123 2714 7123 0 chanx_left_in[19]
rlabel via1 2898 2482 2898 2482 0 chanx_left_in[1]
rlabel metal1 2185 5678 2185 5678 0 chanx_left_in[20]
rlabel metal1 3358 6426 3358 6426 0 chanx_left_in[21]
rlabel metal3 2062 10540 2062 10540 0 chanx_left_in[22]
rlabel metal3 828 10880 828 10880 0 chanx_left_in[23]
rlabel metal3 1717 11356 1717 11356 0 chanx_left_in[24]
rlabel metal1 3082 5644 3082 5644 0 chanx_left_in[25]
rlabel metal2 1794 10557 1794 10557 0 chanx_left_in[26]
rlabel metal3 1717 12580 1717 12580 0 chanx_left_in[27]
rlabel metal2 3266 12920 3266 12920 0 chanx_left_in[28]
rlabel metal1 1380 12818 1380 12818 0 chanx_left_in[29]
rlabel metal1 1610 2550 1610 2550 0 chanx_left_in[2]
rlabel metal1 1610 2924 1610 2924 0 chanx_left_in[3]
rlabel metal1 4140 3502 4140 3502 0 chanx_left_in[4]
rlabel metal3 1004 3604 1004 3604 0 chanx_left_in[5]
rlabel metal2 1242 3553 1242 3553 0 chanx_left_in[6]
rlabel metal2 3726 4267 3726 4267 0 chanx_left_in[7]
rlabel metal2 1610 4471 1610 4471 0 chanx_left_in[8]
rlabel metal3 1004 5236 1004 5236 0 chanx_left_in[9]
rlabel metal3 1372 13804 1372 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal2 2806 18819 2806 18819 0 chanx_left_out[11]
rlabel metal2 2898 19227 2898 19227 0 chanx_left_out[12]
rlabel metal3 1694 19108 1694 19108 0 chanx_left_out[13]
rlabel metal2 2990 19703 2990 19703 0 chanx_left_out[14]
rlabel metal2 3358 20689 3358 20689 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 3726 22015 3726 22015 0 chanx_left_out[20]
rlabel metal1 4002 20978 4002 20978 0 chanx_left_out[21]
rlabel metal1 6854 20366 6854 20366 0 chanx_left_out[22]
rlabel metal1 3910 21114 3910 21114 0 chanx_left_out[23]
rlabel metal1 7544 19890 7544 19890 0 chanx_left_out[24]
rlabel metal1 4324 17238 4324 17238 0 chanx_left_out[25]
rlabel metal1 4830 16558 4830 16558 0 chanx_left_out[26]
rlabel metal1 5474 17714 5474 17714 0 chanx_left_out[27]
rlabel metal2 3174 25041 3174 25041 0 chanx_left_out[28]
rlabel metal1 9890 20842 9890 20842 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 912 15028 912 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal2 22172 18836 22172 18836 0 chany_top_in[0]
rlabel metal1 36432 21590 36432 21590 0 chany_top_in[10]
rlabel metal2 36938 24208 36938 24208 0 chany_top_in[11]
rlabel metal1 32430 21590 32430 21590 0 chany_top_in[12]
rlabel metal2 42458 23970 42458 23970 0 chany_top_in[13]
rlabel metal1 38042 23698 38042 23698 0 chany_top_in[14]
rlabel metal2 37398 21597 37398 21597 0 chany_top_in[15]
rlabel metal1 34408 22202 34408 22202 0 chany_top_in[16]
rlabel metal1 34822 24106 34822 24106 0 chany_top_in[17]
rlabel metal1 37168 21658 37168 21658 0 chany_top_in[18]
rlabel metal1 35687 23698 35687 23698 0 chany_top_in[19]
rlabel metal2 32246 24174 32246 24174 0 chany_top_in[1]
rlabel metal1 37490 24106 37490 24106 0 chany_top_in[20]
rlabel metal1 39882 22474 39882 22474 0 chany_top_in[21]
rlabel metal1 36616 21522 36616 21522 0 chany_top_in[22]
rlabel metal1 40986 23120 40986 23120 0 chany_top_in[23]
rlabel metal1 38180 21998 38180 21998 0 chany_top_in[24]
rlabel metal1 38410 24174 38410 24174 0 chany_top_in[25]
rlabel metal1 39100 24174 39100 24174 0 chany_top_in[26]
rlabel metal1 40158 23630 40158 23630 0 chany_top_in[27]
rlabel metal1 40802 24174 40802 24174 0 chany_top_in[28]
rlabel metal1 42182 23120 42182 23120 0 chany_top_in[29]
rlabel via2 1610 11101 1610 11101 0 chany_top_in[2]
rlabel metal3 12788 7208 12788 7208 0 chany_top_in[3]
rlabel metal1 39790 22066 39790 22066 0 chany_top_in[4]
rlabel metal2 25438 24881 25438 24881 0 chany_top_in[5]
rlabel metal3 16284 23120 16284 23120 0 chany_top_in[6]
rlabel metal2 35098 23732 35098 23732 0 chany_top_in[7]
rlabel metal2 29118 24446 29118 24446 0 chany_top_in[8]
rlabel metal1 36386 24174 36386 24174 0 chany_top_in[9]
rlabel metal1 3772 21454 3772 21454 0 chany_top_out[0]
rlabel metal1 8786 24242 8786 24242 0 chany_top_out[10]
rlabel metal1 9568 23766 9568 23766 0 chany_top_out[11]
rlabel metal2 10718 24497 10718 24497 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal1 12190 20978 12190 20978 0 chany_top_out[14]
rlabel metal2 12558 25034 12558 25034 0 chany_top_out[15]
rlabel metal2 13301 26316 13301 26316 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13984 24242 13984 24242 0 chany_top_out[18]
rlabel metal1 15410 22134 15410 22134 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal1 17342 20978 17342 20978 0 chany_top_out[22]
rlabel metal1 16928 23018 16928 23018 0 chany_top_out[23]
rlabel metal1 16238 23630 16238 23630 0 chany_top_out[24]
rlabel metal1 16192 24106 16192 24106 0 chany_top_out[25]
rlabel metal1 18676 23766 18676 23766 0 chany_top_out[26]
rlabel metal1 20700 22066 20700 22066 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 21574 25272 21574 25272 0 chany_top_out[29]
rlabel metal1 4094 23698 4094 23698 0 chany_top_out[2]
rlabel metal1 5428 22678 5428 22678 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7130 22134 7130 22134 0 chany_top_out[6]
rlabel metal1 6348 24242 6348 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8694 24422 8694 24422 0 chany_top_out[9]
rlabel metal1 17204 21318 17204 21318 0 clknet_0_prog_clk
rlabel metal2 8418 6256 8418 6256 0 clknet_4_0_0_prog_clk
rlabel metal1 24932 14926 24932 14926 0 clknet_4_10_0_prog_clk
rlabel metal2 21114 16082 21114 16082 0 clknet_4_11_0_prog_clk
rlabel metal1 16284 17714 16284 17714 0 clknet_4_12_0_prog_clk
rlabel metal1 20700 18802 20700 18802 0 clknet_4_13_0_prog_clk
rlabel metal1 28244 20434 28244 20434 0 clknet_4_14_0_prog_clk
rlabel metal1 38134 21658 38134 21658 0 clknet_4_15_0_prog_clk
rlabel metal2 9338 13056 9338 13056 0 clknet_4_1_0_prog_clk
rlabel metal1 17112 11118 17112 11118 0 clknet_4_2_0_prog_clk
rlabel metal1 14720 13362 14720 13362 0 clknet_4_3_0_prog_clk
rlabel metal1 6578 18122 6578 18122 0 clknet_4_4_0_prog_clk
rlabel metal1 8602 20298 8602 20298 0 clknet_4_5_0_prog_clk
rlabel metal1 14628 18190 14628 18190 0 clknet_4_6_0_prog_clk
rlabel metal1 13202 21590 13202 21590 0 clknet_4_7_0_prog_clk
rlabel metal1 20792 11118 20792 11118 0 clknet_4_8_0_prog_clk
rlabel metal2 20286 13090 20286 13090 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 2414 25576 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28382 1581 28382 1581 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 2414 33580 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal1 14812 5746 14812 5746 0 gfpga_pad_io_soc_out[0]
rlabel metal2 17434 2710 17434 2710 0 gfpga_pad_io_soc_out[1]
rlabel metal1 19412 4046 19412 4046 0 gfpga_pad_io_soc_out[2]
rlabel metal1 21574 2958 21574 2958 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal1 4278 2312 4278 2312 0 net1
rlabel metal2 9706 17408 9706 17408 0 net10
rlabel metal1 17250 18870 17250 18870 0 net100
rlabel metal1 12696 19754 12696 19754 0 net101
rlabel metal2 3450 15215 3450 15215 0 net102
rlabel metal2 3542 14756 3542 14756 0 net103
rlabel metal2 3358 16354 3358 16354 0 net104
rlabel metal2 13846 16745 13846 16745 0 net105
rlabel metal2 1794 18326 1794 18326 0 net106
rlabel metal1 2277 17646 2277 17646 0 net107
rlabel metal1 1794 18292 1794 18292 0 net108
rlabel metal2 2346 14994 2346 14994 0 net109
rlabel metal2 13386 15861 13386 15861 0 net11
rlabel metal4 16652 15572 16652 15572 0 net110
rlabel metal2 36570 15181 36570 15181 0 net111
rlabel metal2 38502 24429 38502 24429 0 net112
rlabel via2 14214 11339 14214 11339 0 net113
rlabel metal4 19780 17272 19780 17272 0 net114
rlabel metal2 32384 20060 32384 20060 0 net115
rlabel metal2 12466 24565 12466 24565 0 net116
rlabel metal3 13639 12988 13639 12988 0 net117
rlabel metal3 14191 16388 14191 16388 0 net118
rlabel metal2 38778 25007 38778 25007 0 net119
rlabel metal1 6716 6630 6716 6630 0 net12
rlabel metal1 2162 9588 2162 9588 0 net120
rlabel metal2 33810 18989 33810 18989 0 net121
rlabel metal1 15548 21862 15548 21862 0 net122
rlabel metal2 506 18667 506 18667 0 net123
rlabel metal1 15502 23120 15502 23120 0 net124
rlabel metal1 35236 22066 35236 22066 0 net125
rlabel metal2 31786 15895 31786 15895 0 net126
rlabel metal1 17342 23698 17342 23698 0 net127
rlabel metal1 14720 20978 14720 20978 0 net128
rlabel metal2 20102 24565 20102 24565 0 net129
rlabel metal2 414 5439 414 5439 0 net13
rlabel metal1 33718 19890 33718 19890 0 net130
rlabel metal2 966 13396 966 13396 0 net131
rlabel metal1 3542 11254 3542 11254 0 net132
rlabel metal2 506 16388 506 16388 0 net133
rlabel metal2 1104 13532 1104 13532 0 net134
rlabel metal2 552 11628 552 11628 0 net135
rlabel metal2 138 10404 138 10404 0 net136
rlabel metal4 1012 13940 1012 13940 0 net137
rlabel metal2 690 14960 690 14960 0 net138
rlabel metal1 4370 2380 4370 2380 0 net139
rlabel metal1 3082 3162 3082 3162 0 net14
rlabel metal1 7682 2414 7682 2414 0 net140
rlabel metal1 9706 2414 9706 2414 0 net141
rlabel metal1 12420 2414 12420 2414 0 net142
rlabel via2 16974 21437 16974 21437 0 net143
rlabel metal1 23552 23630 23552 23630 0 net144
rlabel metal4 1196 13668 1196 13668 0 net145
rlabel metal1 21298 22644 21298 22644 0 net146
rlabel metal1 21574 24038 21574 24038 0 net147
rlabel metal1 21666 22984 21666 22984 0 net148
rlabel metal1 25530 21658 25530 21658 0 net149
rlabel metal2 1886 5916 1886 5916 0 net15
rlabel metal1 31993 20978 31993 20978 0 net150
rlabel metal1 27462 18394 27462 18394 0 net151
rlabel metal1 18906 13158 18906 13158 0 net152
rlabel metal2 21298 17748 21298 17748 0 net153
rlabel metal1 24334 18802 24334 18802 0 net154
rlabel metal1 13294 20502 13294 20502 0 net155
rlabel metal1 20010 14042 20010 14042 0 net156
rlabel metal2 14306 7616 14306 7616 0 net157
rlabel metal1 14490 6426 14490 6426 0 net158
rlabel metal1 10120 6426 10120 6426 0 net159
rlabel metal2 9890 16915 9890 16915 0 net16
rlabel metal2 10718 6698 10718 6698 0 net160
rlabel metal1 20838 12886 20838 12886 0 net161
rlabel metal1 14858 7854 14858 7854 0 net162
rlabel metal1 16606 13362 16606 13362 0 net163
rlabel metal1 15594 16490 15594 16490 0 net164
rlabel metal1 8280 16218 8280 16218 0 net165
rlabel metal1 10212 7514 10212 7514 0 net166
rlabel metal1 9476 13158 9476 13158 0 net167
rlabel metal1 11776 15334 11776 15334 0 net168
rlabel metal1 10718 6290 10718 6290 0 net169
rlabel metal1 6164 16218 6164 16218 0 net17
rlabel metal1 5888 8602 5888 8602 0 net170
rlabel metal2 14030 8874 14030 8874 0 net171
rlabel metal1 736 10642 736 10642 0 net172
rlabel metal1 11822 6426 11822 6426 0 net173
rlabel metal2 15778 17204 15778 17204 0 net174
rlabel metal1 36110 21658 36110 21658 0 net175
rlabel metal2 10166 19295 10166 19295 0 net176
rlabel metal1 10856 17510 10856 17510 0 net177
rlabel metal1 8418 12308 8418 12308 0 net178
rlabel metal2 12466 13464 12466 13464 0 net179
rlabel metal1 2070 7378 2070 7378 0 net18
rlabel metal1 20562 12750 20562 12750 0 net180
rlabel metal1 16008 7446 16008 7446 0 net181
rlabel metal2 7222 9350 7222 9350 0 net182
rlabel metal1 5934 13158 5934 13158 0 net183
rlabel metal1 14536 17170 14536 17170 0 net184
rlabel metal2 15686 19227 15686 19227 0 net185
rlabel metal1 28060 16558 28060 16558 0 net186
rlabel metal3 14260 20740 14260 20740 0 net187
rlabel metal1 2346 7922 2346 7922 0 net188
rlabel metal1 18814 19482 18814 19482 0 net189
rlabel metal1 1932 6834 1932 6834 0 net19
rlabel metal2 18998 15810 18998 15810 0 net190
rlabel metal1 33442 24038 33442 24038 0 net191
rlabel metal2 26266 21352 26266 21352 0 net192
rlabel metal1 23046 18190 23046 18190 0 net193
rlabel metal1 13110 10574 13110 10574 0 net194
rlabel metal1 32936 24378 32936 24378 0 net195
rlabel metal3 11155 13668 11155 13668 0 net196
rlabel metal1 15180 14450 15180 14450 0 net197
rlabel metal2 22586 7072 22586 7072 0 net198
rlabel metal2 32154 20213 32154 20213 0 net199
rlabel metal2 48714 23018 48714 23018 0 net2
rlabel metal2 2714 11356 2714 11356 0 net20
rlabel metal1 26082 14926 26082 14926 0 net200
rlabel metal1 8050 12750 8050 12750 0 net201
rlabel via2 1610 24293 1610 24293 0 net202
rlabel metal2 3450 11560 3450 11560 0 net203
rlabel metal1 10258 15980 10258 15980 0 net204
rlabel metal1 15640 4794 15640 4794 0 net205
rlabel metal3 8809 19380 8809 19380 0 net206
rlabel metal3 6371 19380 6371 19380 0 net207
rlabel metal1 33120 21862 33120 21862 0 net208
rlabel metal2 22586 14552 22586 14552 0 net209
rlabel metal1 1518 10098 1518 10098 0 net21
rlabel metal2 20010 18972 20010 18972 0 net210
rlabel metal1 14076 15062 14076 15062 0 net211
rlabel metal1 5382 10234 5382 10234 0 net212
rlabel metal2 18906 19465 18906 19465 0 net213
rlabel metal1 17204 22678 17204 22678 0 net214
rlabel metal1 12006 13226 12006 13226 0 net215
rlabel metal1 22126 17578 22126 17578 0 net216
rlabel metal1 22724 10778 22724 10778 0 net217
rlabel metal1 28750 20536 28750 20536 0 net218
rlabel metal1 27225 18938 27225 18938 0 net219
rlabel metal1 4370 15470 4370 15470 0 net22
rlabel metal2 7498 14144 7498 14144 0 net220
rlabel metal3 5290 15844 5290 15844 0 net221
rlabel metal1 16422 8602 16422 8602 0 net222
rlabel metal2 12558 20196 12558 20196 0 net223
rlabel metal1 2392 12410 2392 12410 0 net224
rlabel metal2 20930 16745 20930 16745 0 net225
rlabel metal2 20010 11492 20010 11492 0 net226
rlabel metal2 3818 13294 3818 13294 0 net227
rlabel metal1 27600 17578 27600 17578 0 net228
rlabel metal2 21482 20060 21482 20060 0 net229
rlabel metal1 2024 8398 2024 8398 0 net23
rlabel metal1 20746 13362 20746 13362 0 net230
rlabel metal3 7429 21012 7429 21012 0 net231
rlabel metal1 13570 8058 13570 8058 0 net232
rlabel metal1 18124 8058 18124 8058 0 net233
rlabel metal1 17250 8602 17250 8602 0 net234
rlabel metal2 12374 6494 12374 6494 0 net235
rlabel metal1 13156 21454 13156 21454 0 net236
rlabel metal1 25070 17578 25070 17578 0 net237
rlabel metal1 19780 16490 19780 16490 0 net238
rlabel metal1 17802 14450 17802 14450 0 net239
rlabel metal1 19596 15606 19596 15606 0 net24
rlabel metal2 17434 15912 17434 15912 0 net240
rlabel metal2 12006 7854 12006 7854 0 net241
rlabel metal2 8602 9316 8602 9316 0 net242
rlabel metal1 23644 21590 23644 21590 0 net243
rlabel metal1 17342 13838 17342 13838 0 net244
rlabel metal1 21114 9146 21114 9146 0 net245
rlabel metal1 28244 23630 28244 23630 0 net246
rlabel metal1 29348 18190 29348 18190 0 net247
rlabel metal2 34730 24004 34730 24004 0 net248
rlabel metal2 33718 22814 33718 22814 0 net249
rlabel metal1 1886 2516 1886 2516 0 net25
rlabel metal2 13432 11186 13432 11186 0 net250
rlabel metal2 17710 20111 17710 20111 0 net251
rlabel metal1 24886 12750 24886 12750 0 net252
rlabel metal1 12052 6834 12052 6834 0 net253
rlabel metal1 15640 7514 15640 7514 0 net254
rlabel metal1 32890 22066 32890 22066 0 net255
rlabel metal1 5106 10778 5106 10778 0 net256
rlabel metal1 5888 18666 5888 18666 0 net257
rlabel metal2 27830 10336 27830 10336 0 net258
rlabel metal1 26811 20026 26811 20026 0 net259
rlabel metal2 14214 9112 14214 9112 0 net26
rlabel metal1 24564 20502 24564 20502 0 net260
rlabel metal1 7544 9146 7544 9146 0 net261
rlabel metal1 34086 21114 34086 21114 0 net262
rlabel metal2 31602 23664 31602 23664 0 net263
rlabel metal2 30498 21658 30498 21658 0 net264
rlabel metal1 28934 19278 28934 19278 0 net265
rlabel metal1 27554 15946 27554 15946 0 net266
rlabel metal1 2392 11866 2392 11866 0 net267
rlabel metal1 26949 22202 26949 22202 0 net268
rlabel metal2 30038 23392 30038 23392 0 net269
rlabel metal1 6992 9894 6992 9894 0 net27
rlabel metal2 33074 23987 33074 23987 0 net270
rlabel via2 20010 22661 20010 22661 0 net271
rlabel metal1 22310 10234 22310 10234 0 net272
rlabel metal2 21390 15266 21390 15266 0 net273
rlabel metal2 22678 20060 22678 20060 0 net274
rlabel metal1 19826 15062 19826 15062 0 net275
rlabel metal2 31694 22695 31694 22695 0 net276
rlabel metal1 14582 23630 14582 23630 0 net277
rlabel metal2 15502 18751 15502 18751 0 net278
rlabel metal1 17158 17238 17158 17238 0 net279
rlabel metal1 1886 3468 1886 3468 0 net28
rlabel metal1 17802 13192 17802 13192 0 net280
rlabel metal2 22678 9860 22678 9860 0 net281
rlabel metal1 8326 9622 8326 9622 0 net282
rlabel metal2 19274 9894 19274 9894 0 net283
rlabel metal1 15824 8058 15824 8058 0 net284
rlabel metal2 3772 19244 3772 19244 0 net285
rlabel metal2 9430 9248 9430 9248 0 net286
rlabel metal1 21988 10574 21988 10574 0 net287
rlabel metal1 24288 11662 24288 11662 0 net288
rlabel metal1 26496 16014 26496 16014 0 net289
rlabel metal1 5336 3162 5336 3162 0 net29
rlabel metal2 13570 7293 13570 7293 0 net3
rlabel metal1 6256 3978 6256 3978 0 net30
rlabel metal1 1978 4114 1978 4114 0 net31
rlabel metal1 1886 4556 1886 4556 0 net32
rlabel metal2 17894 21369 17894 21369 0 net33
rlabel metal3 13133 10948 13133 10948 0 net34
rlabel metal1 19734 18156 19734 18156 0 net35
rlabel metal1 8556 21930 8556 21930 0 net36
rlabel metal2 40066 24684 40066 24684 0 net37
rlabel metal1 36892 23562 36892 23562 0 net38
rlabel metal1 36892 23222 36892 23222 0 net39
rlabel metal1 1886 5270 1886 5270 0 net4
rlabel metal1 32706 22032 32706 22032 0 net40
rlabel metal1 12788 12954 12788 12954 0 net41
rlabel metal2 36570 24786 36570 24786 0 net42
rlabel metal2 35926 24616 35926 24616 0 net43
rlabel metal1 23000 20978 23000 20978 0 net44
rlabel metal1 33534 22440 33534 22440 0 net45
rlabel metal2 37306 22865 37306 22865 0 net46
rlabel metal1 34960 21386 34960 21386 0 net47
rlabel metal1 32246 20366 32246 20366 0 net48
rlabel metal1 37720 21862 37720 21862 0 net49
rlabel metal1 1886 6324 1886 6324 0 net5
rlabel metal2 12466 19771 12466 19771 0 net50
rlabel metal1 16192 19346 16192 19346 0 net51
rlabel metal1 18722 21896 18722 21896 0 net52
rlabel metal2 41538 18513 41538 18513 0 net53
rlabel metal2 41998 21352 41998 21352 0 net54
rlabel metal2 1886 11407 1886 11407 0 net55
rlabel metal2 16054 21284 16054 21284 0 net56
rlabel metal1 39974 22950 39974 22950 0 net57
rlabel metal1 28750 23800 28750 23800 0 net58
rlabel metal2 14306 24548 14306 24548 0 net59
rlabel metal1 6992 4726 6992 4726 0 net6
rlabel metal2 32798 22831 32798 22831 0 net60
rlabel metal1 25806 22508 25806 22508 0 net61
rlabel metal1 14490 23086 14490 23086 0 net62
rlabel metal1 25162 5066 25162 5066 0 net63
rlabel metal1 27876 2618 27876 2618 0 net64
rlabel metal1 29992 2618 29992 2618 0 net65
rlabel metal1 33212 2618 33212 2618 0 net66
rlabel metal1 32568 2482 32568 2482 0 net67
rlabel metal2 43930 23358 43930 23358 0 net68
rlabel metal1 45356 24038 45356 24038 0 net69
rlabel metal1 7176 5882 7176 5882 0 net7
rlabel metal2 42550 21386 42550 21386 0 net70
rlabel metal2 43562 20230 43562 20230 0 net71
rlabel metal2 46966 19720 46966 19720 0 net72
rlabel metal2 47058 20774 47058 20774 0 net73
rlabel metal1 48668 24038 48668 24038 0 net74
rlabel metal2 43746 21046 43746 21046 0 net75
rlabel metal1 43976 23562 43976 23562 0 net76
rlabel metal1 47794 21522 47794 21522 0 net77
rlabel metal1 5980 18190 5980 18190 0 net78
rlabel metal2 1794 13345 1794 13345 0 net79
rlabel metal2 6486 14722 6486 14722 0 net8
rlabel metal1 1840 18734 1840 18734 0 net80
rlabel metal1 1794 19380 1794 19380 0 net81
rlabel metal1 2162 19822 2162 19822 0 net82
rlabel metal1 1886 20434 1886 20434 0 net83
rlabel metal2 4186 20434 4186 20434 0 net84
rlabel metal1 1794 21556 1794 21556 0 net85
rlabel metal2 6210 21182 6210 21182 0 net86
rlabel metal1 1794 21964 1794 21964 0 net87
rlabel metal1 2622 22610 2622 22610 0 net88
rlabel metal1 2277 23086 2277 23086 0 net89
rlabel metal1 6118 6086 6118 6086 0 net9
rlabel metal2 12834 13515 12834 13515 0 net90
rlabel metal1 16974 19142 16974 19142 0 net91
rlabel metal1 4094 11322 4094 11322 0 net92
rlabel metal1 2484 10710 2484 10710 0 net93
rlabel metal2 21390 24174 21390 24174 0 net94
rlabel metal1 13846 20264 13846 20264 0 net95
rlabel metal1 4600 17170 4600 17170 0 net96
rlabel metal1 4094 16524 4094 16524 0 net97
rlabel metal2 14674 19737 14674 19737 0 net98
rlabel metal2 10534 15232 10534 15232 0 net99
rlabel metal2 38778 2098 38778 2098 0 prog_clk
rlabel metal1 42136 24174 42136 24174 0 prog_reset
rlabel metal2 19642 17884 19642 17884 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 22034 18156 22034 18156 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 29486 16626 29486 16626 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal2 18906 21913 18906 21913 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal2 1702 9214 1702 9214 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 2162 23766 2162 23766 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel via2 19826 23477 19826 23477 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel via2 31970 21947 31970 21947 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 20102 20026 20102 20026 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal2 21482 22304 21482 22304 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal2 19182 21641 19182 21641 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal1 33442 24140 33442 24140 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 23920 21454 23920 21454 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 22034 22678 22034 22678 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 26680 18802 26680 18802 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 27738 20434 27738 20434 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel via2 21942 20043 21942 20043 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 21666 20434 21666 20434 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 27646 21114 27646 21114 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal2 27830 20740 27830 20740 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal2 26634 24174 26634 24174 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal2 31970 22644 31970 22644 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal1 32338 23732 32338 23732 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal2 31142 23018 31142 23018 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 30682 21998 30682 21998 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 33074 23052 33074 23052 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 29762 20944 29762 20944 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal1 31234 21420 31234 21420 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 29072 18802 29072 18802 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 31096 18734 31096 18734 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 17296 20366 17296 20366 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel via2 32338 21539 32338 21539 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 29900 17850 29900 17850 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal1 20102 18632 20102 18632 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 21160 19482 21160 19482 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 16146 21420 16146 21420 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 25484 15878 25484 15878 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal2 32430 19074 32430 19074 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal2 27186 15776 27186 15776 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20838 13804 20838 13804 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17756 10438 17756 10438 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal2 23874 14450 23874 14450 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 17066 10574 17066 10574 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 16698 8466 16698 8466 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 20700 14450 20700 14450 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 15870 9486 15870 9486 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal1 16100 7854 16100 7854 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 16376 11322 16376 11322 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal1 19688 14450 19688 14450 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 18354 16014 18354 16014 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 18308 8942 18308 8942 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 20838 8942 20838 8942 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 25714 13804 25714 13804 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 22034 9044 22034 9044 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal2 17802 16116 17802 16116 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal1 16836 15538 16836 15538 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 16008 16626 16008 16626 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 15548 15538 15548 15538 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15594 13498 15594 13498 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal2 7774 14620 7774 14620 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal2 12742 10421 12742 10421 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal1 13662 9010 13662 9010 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 12236 10778 12236 10778 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal1 12972 9894 12972 9894 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 13708 13430 13708 13430 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 13616 11186 13616 11186 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 3634 12699 3634 12699 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal1 8602 15096 8602 15096 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 11500 7854 11500 7854 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 14076 16150 14076 16150 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 9936 20366 9936 20366 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal1 12052 19686 12052 19686 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel via2 7314 18581 7314 18581 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 9016 19482 9016 19482 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 16422 12750 16422 12750 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 22586 13804 22586 13804 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 17664 12750 17664 12750 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 7360 21386 7360 21386 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal1 8418 16660 8418 16660 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal3 17204 23800 17204 23800 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel via2 12558 21573 12558 21573 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal3 12834 21352 12834 21352 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 16330 19414 16330 19414 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 1748 9622 1748 9622 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14168 20502 14168 20502 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 17204 18598 17204 18598 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal1 19412 17646 19412 17646 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal2 20470 17918 20470 17918 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 21252 14926 21252 14926 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal2 23966 15164 23966 15164 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 19044 16082 19044 16082 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 25760 15538 25760 15538 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal2 21758 9554 21758 9554 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal2 10534 16949 10534 16949 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 26358 19686 26358 19686 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27922 16422 27922 16422 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21597 19686 21597 19686 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16054 20383 16054 20383 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 19550 23392 19550 23392 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35604 20570 35604 20570 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15410 24378 15410 24378 0 sb_8__0_.mux_left_track_13.out
rlabel metal1 15134 20978 15134 20978 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14766 20825 14766 20825 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2024 10642 2024 10642 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 19366 19822 19366 19822 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 32430 19669 32430 19669 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4968 9146 4968 9146 0 sb_8__0_.mux_left_track_17.out
rlabel metal1 20010 22406 20010 22406 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 18469 18020 18469 18020 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17158 19346 17158 19346 0 sb_8__0_.mux_left_track_19.out
rlabel metal1 23736 21658 23736 21658 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 16082 21528 16082 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11960 7514 11960 7514 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 23414 19482 23414 19482 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 12788 6936 12788 6936 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 12926 13821 12926 13821 0 sb_8__0_.mux_left_track_3.out
rlabel metal1 16422 21012 16422 21012 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16422 19261 16422 19261 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 15334 7866 15334 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 24426 19822 24426 19822 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22724 13940 22724 13940 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4002 5848 4002 5848 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 24012 21998 24012 21998 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4186 5729 4186 5729 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4048 6426 4048 6426 0 sb_8__0_.mux_left_track_35.out
rlabel metal1 30498 22474 30498 22474 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 4186 6307 4186 6307 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 13938 14875 13938 14875 0 sb_8__0_.mux_left_track_45.out
rlabel metal2 30038 21760 30038 21760 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14122 15079 14122 15079 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13754 17272 13754 17272 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 25208 20978 25208 20978 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 17340 24610 17340 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5152 13226 5152 13226 0 sb_8__0_.mux_left_track_49.out
rlabel metal1 29026 18666 29026 18666 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 12342 19458 12342 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 4370 15317 4370 15317 0 sb_8__0_.mux_left_track_5.out
rlabel metal2 17526 20944 17526 20944 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 17135 19380 17135 19380 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5980 13294 5980 13294 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 26496 17306 26496 17306 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 14076 14960 14076 14960 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8418 17918 8418 17918 0 sb_8__0_.mux_left_track_7.out
rlabel metal2 18630 18734 18630 18734 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 18538 18938 18538 18938 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14950 18734 14950 18734 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9154 21454 9154 21454 0 sb_8__0_.mux_left_track_9.out
rlabel metal1 14306 20570 14306 20570 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12650 20230 12650 20230 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31694 19975 31694 19975 0 sb_8__0_.mux_top_track_0.out
rlabel metal1 27738 16660 27738 16660 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28520 16490 28520 16490 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25714 16218 25714 16218 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21091 16218 21091 16218 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23230 15946 23230 15946 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 34822 21930 34822 21930 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 18906 12682 18906 12682 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23322 13056 23322 13056 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16652 10710 16652 10710 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15226 10710 15226 10710 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15778 10506 15778 10506 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel via2 32890 23851 32890 23851 0 sb_8__0_.mux_top_track_12.out
rlabel metal3 16790 12580 16790 12580 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14536 8058 14536 8058 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13846 10778 13846 10778 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13570 10370 13570 10370 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 16008 11594 16008 11594 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10258 9724 10258 9724 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29670 16558 29670 16558 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 34776 21522 34776 21522 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 13938 12206 13938 12206 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 11322 12926 11322 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12880 9010 12880 9010 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33718 17187 33718 17187 0 sb_8__0_.mux_top_track_18.out
rlabel metal1 18492 16218 18492 16218 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14260 13770 14260 13770 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13570 14246 13570 14246 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 1518 9605 1518 9605 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 25438 13158 25438 13158 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25024 13294 25024 13294 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 9588 21022 9588 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13524 8330 13524 8330 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26036 16626 26036 16626 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal3 12604 7344 12604 7344 0 sb_8__0_.mux_top_track_20.out
rlabel metal2 15962 16388 15962 16388 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16744 16966 16744 16966 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel via1 35650 20366 35650 20366 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 15134 15674 15134 15674 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel via3 15019 15300 15019 15300 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35650 20298 35650 20298 0 sb_8__0_.mux_top_track_24.out
rlabel metal1 15364 14042 15364 14042 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18446 11764 18446 11764 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37214 21386 37214 21386 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 10442 11730 10442 11730 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7774 8466 7774 8466 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35604 20842 35604 20842 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 9890 13158 9890 13158 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9200 13158 9200 13158 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 37582 21250 37582 21250 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12466 11849 12466 11849 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12190 15385 12190 15385 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 38962 21165 38962 21165 0 sb_8__0_.mux_top_track_32.out
rlabel metal2 12282 15351 12282 15351 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 28658 18921 28658 18921 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37950 22202 37950 22202 0 sb_8__0_.mux_top_track_34.out
rlabel metal2 12466 17255 12466 17255 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37950 21318 37950 21318 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36708 20842 36708 20842 0 sb_8__0_.mux_top_track_36.out
rlabel metal2 9752 17884 9752 17884 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 6003 18020 6003 18020 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 7682 7412 7682 7412 0 sb_8__0_.mux_top_track_38.out
rlabel metal2 8510 18802 8510 18802 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 1196 16932 1196 16932 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel via3 13547 15300 13547 15300 0 sb_8__0_.mux_top_track_4.out
rlabel metal2 17618 13226 17618 13226 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17526 13311 17526 13311 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16606 12954 16606 12954 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15732 12818 15732 12818 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 15594 14212 15594 14212 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5382 6630 5382 6630 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7774 16422 7774 16422 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21942 8041 21942 8041 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1886 8058 1886 8058 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 11500 21658 11500 21658 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1564 7854 1564 7854 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 37076 21964 37076 21964 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 15962 19482 15962 19482 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9798 20502 9798 20502 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 37122 17017 37122 17017 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33304 19142 33304 19142 0 sb_8__0_.mux_top_track_46.out
rlabel metal1 17342 18054 17342 18054 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10580 17510 10580 17510 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13018 19737 13018 19737 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5566 9044 5566 9044 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 19550 18394 19550 18394 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12098 16694 12098 16694 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15732 18054 15732 18054 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 35098 15385 35098 15385 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 20746 17578 20746 17578 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14996 16694 14996 16694 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 16882 18139 16882 18139 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40112 23698 40112 23698 0 sb_8__0_.mux_top_track_6.out
rlabel metal1 23092 16082 23092 16082 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22908 16218 22908 16218 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20194 15742 20194 15742 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14812 12954 14812 12954 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19504 15334 19504 15334 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 29670 16949 29670 16949 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 24932 12274 24932 12274 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel via1 24978 12189 24978 12189 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21367 13906 21367 13906 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14674 9078 14674 9078 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20194 13804 20194 13804 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 44758 25340 44758 25340 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45494 25296 45494 25296 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46368 24174 46368 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 46736 23698 46736 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48254 24174 48254 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 43378 23834 43378 23834 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44252 23698 44252 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 46874 21437 46874 21437 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 45494 20315 45494 20315 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 47357 23732 47357 23732 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 45862 22015 45862 22015 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2234 41446 2234 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2200 44114 2200 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 46782 2166 46782 2166 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49450 2132 49450 2132 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
